// author Mace

module SNAX_DIMC # (
    parameter int unsigned NarrowDataWidth = 64,
    parameter int unsigned WideDataWidth   = 512,
    parameter int unsigned RegAddrWidth    = 32,
    parameter int unsigned RegDataWidth    = 32
)(
    clk_i, rst_ni,
    acc2stream_0_data_o, acc2stream_0_valid_o, acc2stream_0_ready_i,
    stream2acc_0_data_i, stream2acc_0_valid_i, stream2acc_0_ready_o,
    stream2acc_1_data_i, stream2acc_1_valid_i, stream2acc_1_ready_o,
    stream2acc_2_data_i, stream2acc_2_valid_i, stream2acc_2_ready_o,
    stream2acc_3_data_i, stream2acc_3_valid_i, stream2acc_3_ready_o,
    csr_req_addr_i, csr_req_data_i, csr_req_write_i, csr_req_valid_i, csr_req_ready_o,
    csr_rsp_data_o, csr_rsp_valid_o, csr_rsp_ready_i
);

/**************************************************************************/
// Clock and reset
/**************************************************************************/
input  logic                       clk_i;
input  logic                       rst_ni;

/**************************************************************************/
// Accelerator ports
/**************************************************************************/
// Ports from accelerator to streamer by writer data movers
output logic [WideDataWidth-1:0]   acc2stream_0_data_o;
output logic                       acc2stream_0_valid_o;
input  logic                       acc2stream_0_ready_i;
    
// Ports from streamer to accelerator by reader data movers
input  logic [WideDataWidth-1:0]   stream2acc_0_data_i;
input  logic                       stream2acc_0_valid_i;
output logic                       stream2acc_0_ready_o;

input  logic [WideDataWidth-1:0]   stream2acc_1_data_i;
input  logic                       stream2acc_1_valid_i;
output logic                       stream2acc_1_ready_o;

input  logic [WideDataWidth-1:0]   stream2acc_2_data_i;
input  logic                       stream2acc_2_valid_i;
output logic                       stream2acc_2_ready_o;

input  logic [WideDataWidth-1:0]   stream2acc_3_data_i;
input  logic                       stream2acc_3_valid_i;
output logic                       stream2acc_3_ready_o;


/**************************************************************************/
// CSR control ports
/**************************************************************************/
// Request
input  logic [   RegAddrWidth-1:0] csr_req_addr_i;
input  logic [   RegDataWidth-1:0] csr_req_data_i;
input  logic                       csr_req_write_i;
input  logic                       csr_req_valid_i;
output logic                       csr_req_ready_o;
// Response
output logic [   RegDataWidth-1:0] csr_rsp_data_o;
output logic                       csr_rsp_valid_o;
input  logic                       csr_rsp_ready_i;
/**************************************************************************/

// Internal signals

wire rst;

assign rst = ~rst_ni;

wire [191:0] result_QKV_0, result_QKV_1, result_QKV_2, result_QKV_3, result_QKV_4, result_QKV_5, result_QKV_6, result_QKV_7, result_QKV_8, result_QKV_9, result_QKV_10, result_QKV_11, result_QKV_12, result_QKV_13, result_QKV_14, result_QKV_15,
             result_QKV_16, result_QKV_17, result_QKV_18, result_QKV_19, result_QKV_20, result_QKV_21, result_QKV_22, result_QKV_23, result_QKV_24, result_QKV_25, result_QKV_26, result_QKV_27, result_QKV_28, result_QKV_29, result_QKV_30, result_QKV_31,
             result_QKT_0, result_QKT_1, result_QKT_2, result_QKT_3;

wire [63:0] WL_QKV_0, WL_QKV_1, WL_QKV_2, WL_QKV_3, WL_QKV_4, WL_QKV_5, WL_QKV_6, WL_QKV_7, WL_QKV_8, WL_QKV_9, WL_QKV_10, WL_QKV_11, WL_QKV_12, WL_QKV_13, WL_QKV_14, WL_QKV_15,
            WL_QKV_16, WL_QKV_17, WL_QKV_18, WL_QKV_19, WL_QKV_20, WL_QKV_21, WL_QKV_22, WL_QKV_23, WL_QKV_24, WL_QKV_25, WL_QKV_26, WL_QKV_27, WL_QKV_28, WL_QKV_29, WL_QKV_30, WL_QKV_31,
            WL_QKT_0, WL_QKT_1, WL_QKT_2, WL_QKT_3;

wire [127:0] wdata_QKV_0, wdata_QKV_1, wdata_QKV_2, wdata_QKV_3, wdata_QKV_4, wdata_QKV_5, wdata_QKV_6, wdata_QKV_7, wdata_QKV_8, wdata_QKV_9, wdata_QKV_10, wdata_QKV_11, wdata_QKV_12, wdata_QKV_13, wdata_QKV_14, wdata_QKV_15,
             wdata_QKV_16, wdata_QKV_17, wdata_QKV_18, wdata_QKV_19, wdata_QKV_20, wdata_QKV_21, wdata_QKV_22, wdata_QKV_23, wdata_QKV_24, wdata_QKV_25, wdata_QKV_26, wdata_QKV_27, wdata_QKV_28, wdata_QKV_29, wdata_QKV_30, wdata_QKV_31,
             wdata_QKT_0, wdata_QKT_1, wdata_QKT_2, wdata_QKT_3;

wire [63:0] ai_QKV_0, ai_QKV_1, ai_QKV_2, ai_QKV_3, ai_QKV_4, ai_QKV_5, ai_QKV_6, ai_QKV_7, ai_QKV_8, ai_QKV_9, ai_QKV_10, ai_QKV_11, ai_QKV_12, ai_QKV_13, ai_QKV_14, ai_QKV_15,
            ai_QKV_16, ai_QKV_17, ai_QKV_18, ai_QKV_19, ai_QKV_20, ai_QKV_21, ai_QKV_22, ai_QKV_23, ai_QKV_24, ai_QKV_25, ai_QKV_26, ai_QKV_27, ai_QKV_28, ai_QKV_29, ai_QKV_30, ai_QKV_31,
            ai_QKT_0, ai_QKT_1, ai_QKT_2, ai_QKT_3;

wire RE_QKV__0, RE_QKV__1, RE_QKV__2, RE_QKV__3, RE_QKV__4, RE_QKV__5, RE_QKV__6, RE_QKV__7, RE_QKV__8, RE_QKV__9, RE_QKV__10, RE_QKV__11, RE_QKV__12, RE_QKV__13, RE_QKV__14, RE_QKV__15,
     RE_QKV__16, RE_QKV__17, RE_QKV__18, RE_QKV__19, RE_QKV__20, RE_QKV__21, RE_QKV__22, RE_QKV__23, RE_QKV__24, RE_QKV__25, RE_QKV__26, RE_QKV__27, RE_QKV__28, RE_QKV__29, RE_QKV__30, RE_QKV__31,
     RE_QKT__0, RE_QKT__1, RE_QKT__2, RE_QKT__3;

wire PREC_QKV_0, PREC_QKV_1, PREC_QKV_2, PREC_QKV_3, PREC_QKV_4, PREC_QKV_5, PREC_QKV_6, PREC_QKV_7, PREC_QKV_8, PREC_QKV_9, PREC_QKV_10, PREC_QKV_11, PREC_QKV_12, PREC_QKV_13, PREC_QKV_14, PREC_QKV_15,
     PREC_QKV_16, PREC_QKV_17, PREC_QKV_18, PREC_QKV_19, PREC_QKV_20, PREC_QKV_21, PREC_QKV_22, PREC_QKV_23, PREC_QKV_24, PREC_QKV_25, PREC_QKV_26, PREC_QKV_27, PREC_QKV_28, PREC_QKV_29, PREC_QKV_30, PREC_QKV_31,
     PREC_QKT_0, PREC_QKT_1, PREC_QKT_2, PREC_QKT_3;

wire PREC_QKV__0, PREC_QKV__1, PREC_QKV__2, PREC_QKV__3, PREC_QKV__4, PREC_QKV__5, PREC_QKV__6, PREC_QKV__7, PREC_QKV__8, PREC_QKV__9, PREC_QKV__10, PREC_QKV__11, PREC_QKV__12, PREC_QKV__13, PREC_QKV__14, PREC_QKV__15,
     PREC_QKV__16, PREC_QKV__17, PREC_QKV__18, PREC_QKV__19, PREC_QKV__20, PREC_QKV__21, PREC_QKV__22, PREC_QKV__23, PREC_QKV__24, PREC_QKV__25, PREC_QKV__26, PREC_QKV__27, PREC_QKV__28, PREC_QKV__29, PREC_QKV__30, PREC_QKV__31,
     PREC_QKT__0, PREC_QKT__1, PREC_QKT__2, PREC_QKT__3;

snax_interfaces i_snax_interfaces(
    .clk(clk_i),
    .rst(rst_ni),

    .snax_acc_req_valid(csr_req_valid_i),
    .snax_acc_req_data_addr(csr_req_addr_i),
    .snax_acc_req_data_wen(csr_req_write_i),
    .snax_acc_req_data_data(csr_req_data_i),
    .snax_acc_req_ready(csr_req_ready_o),

    .acc_snax_rsp_valid(csr_rsp_valid_o),
    .acc_snax_rsp_data_data(csr_rsp_data_o),
    .acc_snax_rsp_ready(csr_rsp_ready_i),

    .stream_acc_port_0_valid(stream2acc_0_valid_i),
    .stream_acc_port_0_data(stream2acc_0_data_i),
    .stream_acc_port_0_ready(stream2acc_0_ready_o),

    .stream_acc_port_1_valid(stream2acc_1_valid_i),
    .stream_acc_port_1_data(stream2acc_1_data_i),
    .stream_acc_port_1_ready(stream2acc_1_ready_o),

    .stream_acc_port_2_valid(stream2acc_2_valid_i),
    .stream_acc_port_2_data(stream2acc_2_data_i),
    .stream_acc_port_2_ready(stream2acc_2_ready_o),

    .stream_acc_port_3_valid(stream2acc_3_valid_i),
    .stream_acc_port_3_data(stream2acc_3_data_i),
    .stream_acc_port_3_ready(stream2acc_3_ready_o),

    .acc_stream_port_valid(acc2stream_0_valid_o),
    .acc_stream_port_data(acc2stream_0_data_o),
    .acc_stream_port_ready(acc2stream_0_ready_i),

    // .result_QKV_0(result_QKV_0), .result_QKV_1(result_QKV_1), .result_QKV_2(result_QKV_2), .result_QKV_3(result_QKV_3), .result_QKV_4(result_QKV_4), .result_QKV_5(result_QKV_5), .result_QKV_6(result_QKV_6), .result_QKV_7(result_QKV_7), .result_QKV_8(result_QKV_8), .result_QKV_9(result_QKV_9), .result_QKV_10(result_QKV_10), .result_QKV_11(result_QKV_11), .result_QKV_12(result_QKV_12), .result_QKV_13(result_QKV_13), .result_QKV_14(result_QKV_14), .result_QKV_15(result_QKV_15),
    // .result_QKV_16(result_QKV_16), .result_QKV_17(result_QKV_17), .result_QKV_18(result_QKV_18), .result_QKV_19(result_QKV_19), .result_QKV_20(result_QKV_20), .result_QKV_21(result_QKV_21), .result_QKV_22(result_QKV_22), .result_QKV_23(result_QKV_23), .result_QKV_24(result_QKV_24), .result_QKV_25(result_QKV_25), .result_QKV_26(result_QKV_26), .result_QKV_27(result_QKV_27), .result_QKV_28(result_QKV_28), .result_QKV_29(result_QKV_29), .result_QKV_30(result_QKV_30), .result_QKV_31(result_QKV_31),
    // .result_QKT_0(result_QKT_0), .result_QKT_1(result_QKT_1), .result_QKT_2(result_QKT_2), .result_QKT_3(result_QKT_3),

    .S0_QKV_0(result_QKV_0[11:0]), .S1_QKV_0(result_QKV_0[23:12]), .S2_QKV_0(result_QKV_0[35:24]), .S3_QKV_0(result_QKV_0[47:36]), .S4_QKV_0(result_QKV_0[59:48]), .S5_QKV_0(result_QKV_0[71:60]), .S6_QKV_0(result_QKV_0[83:72]), .S7_QKV_0(result_QKV_0[95:84]), .S8_QKV_0(result_QKV_0[107:96]), .S9_QKV_0(result_QKV_0[119:108]), .S10_QKV_0(result_QKV_0[131:120]), .S11_QKV_0(result_QKV_0[143:132]), .S12_QKV_0(result_QKV_0[155:144]), .S13_QKV_0(result_QKV_0[167:156]), .S14_QKV_0(result_QKV_0[179:168]), .S15_QKV_0(result_QKV_0[191:180]),
    .S0_QKV_1(result_QKV_1[11:0]), .S1_QKV_1(result_QKV_1[23:12]), .S2_QKV_1(result_QKV_1[35:24]), .S3_QKV_1(result_QKV_1[47:36]), .S4_QKV_1(result_QKV_1[59:48]), .S5_QKV_1(result_QKV_1[71:60]), .S6_QKV_1(result_QKV_1[83:72]), .S7_QKV_1(result_QKV_1[95:84]), .S8_QKV_1(result_QKV_1[107:96]), .S9_QKV_1(result_QKV_1[119:108]), .S10_QKV_1(result_QKV_1[131:120]), .S11_QKV_1(result_QKV_1[143:132]), .S12_QKV_1(result_QKV_1[155:144]), .S13_QKV_1(result_QKV_1[167:156]), .S14_QKV_1(result_QKV_1[179:168]), .S15_QKV_1(result_QKV_1[191:180]),
    .S0_QKV_2(result_QKV_2[11:0]), .S1_QKV_2(result_QKV_2[23:12]), .S2_QKV_2(result_QKV_2[35:24]), .S3_QKV_2(result_QKV_2[47:36]), .S4_QKV_2(result_QKV_2[59:48]), .S5_QKV_2(result_QKV_2[71:60]), .S6_QKV_2(result_QKV_2[83:72]), .S7_QKV_2(result_QKV_2[95:84]), .S8_QKV_2(result_QKV_2[107:96]), .S9_QKV_2(result_QKV_2[119:108]), .S10_QKV_2(result_QKV_2[131:120]), .S11_QKV_2(result_QKV_2[143:132]), .S12_QKV_2(result_QKV_2[155:144]), .S13_QKV_2(result_QKV_2[167:156]), .S14_QKV_2(result_QKV_2[179:168]), .S15_QKV_2(result_QKV_2[191:180]),
    .S0_QKV_3(result_QKV_3[11:0]), .S1_QKV_3(result_QKV_3[23:12]), .S2_QKV_3(result_QKV_3[35:24]), .S3_QKV_3(result_QKV_3[47:36]), .S4_QKV_3(result_QKV_3[59:48]), .S5_QKV_3(result_QKV_3[71:60]), .S6_QKV_3(result_QKV_3[83:72]), .S7_QKV_3(result_QKV_3[95:84]), .S8_QKV_3(result_QKV_3[107:96]), .S9_QKV_3(result_QKV_3[119:108]), .S10_QKV_3(result_QKV_3[131:120]), .S11_QKV_3(result_QKV_3[143:132]), .S12_QKV_3(result_QKV_3[155:144]), .S13_QKV_3(result_QKV_3[167:156]), .S14_QKV_3(result_QKV_3[179:168]), .S15_QKV_3(result_QKV_3[191:180]),
    .S0_QKV_4(result_QKV_4[11:0]), .S1_QKV_4(result_QKV_4[23:12]), .S2_QKV_4(result_QKV_4[35:24]), .S3_QKV_4(result_QKV_4[47:36]), .S4_QKV_4(result_QKV_4[59:48]), .S5_QKV_4(result_QKV_4[71:60]), .S6_QKV_4(result_QKV_4[83:72]), .S7_QKV_4(result_QKV_4[95:84]), .S8_QKV_4(result_QKV_4[107:96]), .S9_QKV_4(result_QKV_4[119:108]), .S10_QKV_4(result_QKV_4[131:120]), .S11_QKV_4(result_QKV_4[143:132]), .S12_QKV_4(result_QKV_4[155:144]), .S13_QKV_4(result_QKV_4[167:156]), .S14_QKV_4(result_QKV_4[179:168]), .S15_QKV_4(result_QKV_4[191:180]),
    .S0_QKV_5(result_QKV_5[11:0]), .S1_QKV_5(result_QKV_5[23:12]), .S2_QKV_5(result_QKV_5[35:24]), .S3_QKV_5(result_QKV_5[47:36]), .S4_QKV_5(result_QKV_5[59:48]), .S5_QKV_5(result_QKV_5[71:60]), .S6_QKV_5(result_QKV_5[83:72]), .S7_QKV_5(result_QKV_5[95:84]), .S8_QKV_5(result_QKV_5[107:96]), .S9_QKV_5(result_QKV_5[119:108]), .S10_QKV_5(result_QKV_5[131:120]), .S11_QKV_5(result_QKV_5[143:132]), .S12_QKV_5(result_QKV_5[155:144]), .S13_QKV_5(result_QKV_5[167:156]), .S14_QKV_5(result_QKV_5[179:168]), .S15_QKV_5(result_QKV_5[191:180]),
    .S0_QKV_6(result_QKV_6[11:0]), .S1_QKV_6(result_QKV_6[23:12]), .S2_QKV_6(result_QKV_6[35:24]), .S3_QKV_6(result_QKV_6[47:36]), .S4_QKV_6(result_QKV_6[59:48]), .S5_QKV_6(result_QKV_6[71:60]), .S6_QKV_6(result_QKV_6[83:72]), .S7_QKV_6(result_QKV_6[95:84]), .S8_QKV_6(result_QKV_6[107:96]), .S9_QKV_6(result_QKV_6[119:108]), .S10_QKV_6(result_QKV_6[131:120]), .S11_QKV_6(result_QKV_6[143:132]), .S12_QKV_6(result_QKV_6[155:144]), .S13_QKV_6(result_QKV_6[167:156]), .S14_QKV_6(result_QKV_6[179:168]), .S15_QKV_6(result_QKV_6[191:180]),
    .S0_QKV_7(result_QKV_7[11:0]), .S1_QKV_7(result_QKV_7[23:12]), .S2_QKV_7(result_QKV_7[35:24]), .S3_QKV_7(result_QKV_7[47:36]), .S4_QKV_7(result_QKV_7[59:48]), .S5_QKV_7(result_QKV_7[71:60]), .S6_QKV_7(result_QKV_7[83:72]), .S7_QKV_7(result_QKV_7[95:84]), .S8_QKV_7(result_QKV_7[107:96]), .S9_QKV_7(result_QKV_7[119:108]), .S10_QKV_7(result_QKV_7[131:120]), .S11_QKV_7(result_QKV_7[143:132]), .S12_QKV_7(result_QKV_7[155:144]), .S13_QKV_7(result_QKV_7[167:156]), .S14_QKV_7(result_QKV_7[179:168]), .S15_QKV_7(result_QKV_7[191:180]),
    .S0_QKV_8(result_QKV_8[11:0]), .S1_QKV_8(result_QKV_8[23:12]), .S2_QKV_8(result_QKV_8[35:24]), .S3_QKV_8(result_QKV_8[47:36]), .S4_QKV_8(result_QKV_8[59:48]), .S5_QKV_8(result_QKV_8[71:60]), .S6_QKV_8(result_QKV_8[83:72]), .S7_QKV_8(result_QKV_8[95:84]), .S8_QKV_8(result_QKV_8[107:96]), .S9_QKV_8(result_QKV_8[119:108]), .S10_QKV_8(result_QKV_8[131:120]), .S11_QKV_8(result_QKV_8[143:132]), .S12_QKV_8(result_QKV_8[155:144]), .S13_QKV_8(result_QKV_8[167:156]), .S14_QKV_8(result_QKV_8[179:168]), .S15_QKV_8(result_QKV_8[191:180]),
    .S0_QKV_9(result_QKV_9[11:0]), .S1_QKV_9(result_QKV_9[23:12]), .S2_QKV_9(result_QKV_9[35:24]), .S3_QKV_9(result_QKV_9[47:36]), .S4_QKV_9(result_QKV_9[59:48]), .S5_QKV_9(result_QKV_9[71:60]), .S6_QKV_9(result_QKV_9[83:72]), .S7_QKV_9(result_QKV_9[95:84]), .S8_QKV_9(result_QKV_9[107:96]), .S9_QKV_9(result_QKV_9[119:108]), .S10_QKV_9(result_QKV_9[131:120]), .S11_QKV_9(result_QKV_9[143:132]), .S12_QKV_9(result_QKV_9[155:144]), .S13_QKV_9(result_QKV_9[167:156]), .S14_QKV_9(result_QKV_9[179:168]), .S15_QKV_9(result_QKV_9[191:180]),
    .S0_QKV_10(result_QKV_10[11:0]), .S1_QKV_10(result_QKV_10[23:12]), .S2_QKV_10(result_QKV_10[35:24]), .S3_QKV_10(result_QKV_10[47:36]), .S4_QKV_10(result_QKV_10[59:48]), .S5_QKV_10(result_QKV_10[71:60]), .S6_QKV_10(result_QKV_10[83:72]), .S7_QKV_10(result_QKV_10[95:84]), .S8_QKV_10(result_QKV_10[107:96]), .S9_QKV_10(result_QKV_10[119:108]), .S10_QKV_10(result_QKV_10[131:120]), .S11_QKV_10(result_QKV_10[143:132]), .S12_QKV_10(result_QKV_10[155:144]), .S13_QKV_10(result_QKV_10[167:156]), .S14_QKV_10(result_QKV_10[179:168]), .S15_QKV_10(result_QKV_10[191:180]),
    .S0_QKV_11(result_QKV_11[11:0]), .S1_QKV_11(result_QKV_11[23:12]), .S2_QKV_11(result_QKV_11[35:24]), .S3_QKV_11(result_QKV_11[47:36]), .S4_QKV_11(result_QKV_11[59:48]), .S5_QKV_11(result_QKV_11[71:60]), .S6_QKV_11(result_QKV_11[83:72]), .S7_QKV_11(result_QKV_11[95:84]), .S8_QKV_11(result_QKV_11[107:96]), .S9_QKV_11(result_QKV_11[119:108]), .S10_QKV_11(result_QKV_11[131:120]), .S11_QKV_11(result_QKV_11[143:132]), .S12_QKV_11(result_QKV_11[155:144]), .S13_QKV_11(result_QKV_11[167:156]), .S14_QKV_11(result_QKV_11[179:168]), .S15_QKV_11(result_QKV_11[191:180]),
    .S0_QKV_12(result_QKV_12[11:0]), .S1_QKV_12(result_QKV_12[23:12]), .S2_QKV_12(result_QKV_12[35:24]), .S3_QKV_12(result_QKV_12[47:36]), .S4_QKV_12(result_QKV_12[59:48]), .S5_QKV_12(result_QKV_12[71:60]), .S6_QKV_12(result_QKV_12[83:72]), .S7_QKV_12(result_QKV_12[95:84]), .S8_QKV_12(result_QKV_12[107:96]), .S9_QKV_12(result_QKV_12[119:108]), .S10_QKV_12(result_QKV_12[131:120]), .S11_QKV_12(result_QKV_12[143:132]), .S12_QKV_12(result_QKV_12[155:144]), .S13_QKV_12(result_QKV_12[167:156]), .S14_QKV_12(result_QKV_12[179:168]), .S15_QKV_12(result_QKV_12[191:180]),
    .S0_QKV_13(result_QKV_13[11:0]), .S1_QKV_13(result_QKV_13[23:12]), .S2_QKV_13(result_QKV_13[35:24]), .S3_QKV_13(result_QKV_13[47:36]), .S4_QKV_13(result_QKV_13[59:48]), .S5_QKV_13(result_QKV_13[71:60]), .S6_QKV_13(result_QKV_13[83:72]), .S7_QKV_13(result_QKV_13[95:84]), .S8_QKV_13(result_QKV_13[107:96]), .S9_QKV_13(result_QKV_13[119:108]), .S10_QKV_13(result_QKV_13[131:120]), .S11_QKV_13(result_QKV_13[143:132]), .S12_QKV_13(result_QKV_13[155:144]), .S13_QKV_13(result_QKV_13[167:156]), .S14_QKV_13(result_QKV_13[179:168]), .S15_QKV_13(result_QKV_13[191:180]),
    .S0_QKV_14(result_QKV_14[11:0]), .S1_QKV_14(result_QKV_14[23:12]), .S2_QKV_14(result_QKV_14[35:24]), .S3_QKV_14(result_QKV_14[47:36]), .S4_QKV_14(result_QKV_14[59:48]), .S5_QKV_14(result_QKV_14[71:60]), .S6_QKV_14(result_QKV_14[83:72]), .S7_QKV_14(result_QKV_14[95:84]), .S8_QKV_14(result_QKV_14[107:96]), .S9_QKV_14(result_QKV_14[119:108]), .S10_QKV_14(result_QKV_14[131:120]), .S11_QKV_14(result_QKV_14[143:132]), .S12_QKV_14(result_QKV_14[155:144]), .S13_QKV_14(result_QKV_14[167:156]), .S14_QKV_14(result_QKV_14[179:168]), .S15_QKV_14(result_QKV_14[191:180]),
    .S0_QKV_15(result_QKV_15[11:0]), .S1_QKV_15(result_QKV_15[23:12]), .S2_QKV_15(result_QKV_15[35:24]), .S3_QKV_15(result_QKV_15[47:36]), .S4_QKV_15(result_QKV_15[59:48]), .S5_QKV_15(result_QKV_15[71:60]), .S6_QKV_15(result_QKV_15[83:72]), .S7_QKV_15(result_QKV_15[95:84]), .S8_QKV_15(result_QKV_15[107:96]), .S9_QKV_15(result_QKV_15[119:108]), .S10_QKV_15(result_QKV_15[131:120]), .S11_QKV_15(result_QKV_15[143:132]), .S12_QKV_15(result_QKV_15[155:144]), .S13_QKV_15(result_QKV_15[167:156]), .S14_QKV_15(result_QKV_15[179:168]), .S15_QKV_15(result_QKV_15[191:180]),
    .S0_QKV_16(result_QKV_16[11:0]), .S1_QKV_16(result_QKV_16[23:12]), .S2_QKV_16(result_QKV_16[35:24]), .S3_QKV_16(result_QKV_16[47:36]), .S4_QKV_16(result_QKV_16[59:48]), .S5_QKV_16(result_QKV_16[71:60]), .S6_QKV_16(result_QKV_16[83:72]), .S7_QKV_16(result_QKV_16[95:84]), .S8_QKV_16(result_QKV_16[107:96]), .S9_QKV_16(result_QKV_16[119:108]), .S10_QKV_16(result_QKV_16[131:120]), .S11_QKV_16(result_QKV_16[143:132]), .S12_QKV_16(result_QKV_16[155:144]), .S13_QKV_16(result_QKV_16[167:156]), .S14_QKV_16(result_QKV_16[179:168]), .S15_QKV_16(result_QKV_16[191:180]),
    .S0_QKV_17(result_QKV_17[11:0]), .S1_QKV_17(result_QKV_17[23:12]), .S2_QKV_17(result_QKV_17[35:24]), .S3_QKV_17(result_QKV_17[47:36]), .S4_QKV_17(result_QKV_17[59:48]), .S5_QKV_17(result_QKV_17[71:60]), .S6_QKV_17(result_QKV_17[83:72]), .S7_QKV_17(result_QKV_17[95:84]), .S8_QKV_17(result_QKV_17[107:96]), .S9_QKV_17(result_QKV_17[119:108]), .S10_QKV_17(result_QKV_17[131:120]), .S11_QKV_17(result_QKV_17[143:132]), .S12_QKV_17(result_QKV_17[155:144]), .S13_QKV_17(result_QKV_17[167:156]), .S14_QKV_17(result_QKV_17[179:168]), .S15_QKV_17(result_QKV_17[191:180]),
    .S0_QKV_18(result_QKV_18[11:0]), .S1_QKV_18(result_QKV_18[23:12]), .S2_QKV_18(result_QKV_18[35:24]), .S3_QKV_18(result_QKV_18[47:36]), .S4_QKV_18(result_QKV_18[59:48]), .S5_QKV_18(result_QKV_18[71:60]), .S6_QKV_18(result_QKV_18[83:72]), .S7_QKV_18(result_QKV_18[95:84]), .S8_QKV_18(result_QKV_18[107:96]), .S9_QKV_18(result_QKV_18[119:108]), .S10_QKV_18(result_QKV_18[131:120]), .S11_QKV_18(result_QKV_18[143:132]), .S12_QKV_18(result_QKV_18[155:144]), .S13_QKV_18(result_QKV_18[167:156]), .S14_QKV_18(result_QKV_18[179:168]), .S15_QKV_18(result_QKV_18[191:180]),
    .S0_QKV_19(result_QKV_19[11:0]), .S1_QKV_19(result_QKV_19[23:12]), .S2_QKV_19(result_QKV_19[35:24]), .S3_QKV_19(result_QKV_19[47:36]), .S4_QKV_19(result_QKV_19[59:48]), .S5_QKV_19(result_QKV_19[71:60]), .S6_QKV_19(result_QKV_19[83:72]), .S7_QKV_19(result_QKV_19[95:84]), .S8_QKV_19(result_QKV_19[107:96]), .S9_QKV_19(result_QKV_19[119:108]), .S10_QKV_19(result_QKV_19[131:120]), .S11_QKV_19(result_QKV_19[143:132]), .S12_QKV_19(result_QKV_19[155:144]), .S13_QKV_19(result_QKV_19[167:156]), .S14_QKV_19(result_QKV_19[179:168]), .S15_QKV_19(result_QKV_19[191:180]),
    .S0_QKV_20(result_QKV_20[11:0]), .S1_QKV_20(result_QKV_20[23:12]), .S2_QKV_20(result_QKV_20[35:24]), .S3_QKV_20(result_QKV_20[47:36]), .S4_QKV_20(result_QKV_20[59:48]), .S5_QKV_20(result_QKV_20[71:60]), .S6_QKV_20(result_QKV_20[83:72]), .S7_QKV_20(result_QKV_20[95:84]), .S8_QKV_20(result_QKV_20[107:96]), .S9_QKV_20(result_QKV_20[119:108]), .S10_QKV_20(result_QKV_20[131:120]), .S11_QKV_20(result_QKV_20[143:132]), .S12_QKV_20(result_QKV_20[155:144]), .S13_QKV_20(result_QKV_20[167:156]), .S14_QKV_20(result_QKV_20[179:168]), .S15_QKV_20(result_QKV_20[191:180]),
    .S0_QKV_21(result_QKV_21[11:0]), .S1_QKV_21(result_QKV_21[23:12]), .S2_QKV_21(result_QKV_21[35:24]), .S3_QKV_21(result_QKV_21[47:36]), .S4_QKV_21(result_QKV_21[59:48]), .S5_QKV_21(result_QKV_21[71:60]), .S6_QKV_21(result_QKV_21[83:72]), .S7_QKV_21(result_QKV_21[95:84]), .S8_QKV_21(result_QKV_21[107:96]), .S9_QKV_21(result_QKV_21[119:108]), .S10_QKV_21(result_QKV_21[131:120]), .S11_QKV_21(result_QKV_21[143:132]), .S12_QKV_21(result_QKV_21[155:144]), .S13_QKV_21(result_QKV_21[167:156]), .S14_QKV_21(result_QKV_21[179:168]), .S15_QKV_21(result_QKV_21[191:180]),
    .S0_QKV_22(result_QKV_22[11:0]), .S1_QKV_22(result_QKV_22[23:12]), .S2_QKV_22(result_QKV_22[35:24]), .S3_QKV_22(result_QKV_22[47:36]), .S4_QKV_22(result_QKV_22[59:48]), .S5_QKV_22(result_QKV_22[71:60]), .S6_QKV_22(result_QKV_22[83:72]), .S7_QKV_22(result_QKV_22[95:84]), .S8_QKV_22(result_QKV_22[107:96]), .S9_QKV_22(result_QKV_22[119:108]), .S10_QKV_22(result_QKV_22[131:120]), .S11_QKV_22(result_QKV_22[143:132]), .S12_QKV_22(result_QKV_22[155:144]), .S13_QKV_22(result_QKV_22[167:156]), .S14_QKV_22(result_QKV_22[179:168]), .S15_QKV_22(result_QKV_22[191:180]),
    .S0_QKV_23(result_QKV_23[11:0]), .S1_QKV_23(result_QKV_23[23:12]), .S2_QKV_23(result_QKV_23[35:24]), .S3_QKV_23(result_QKV_23[47:36]), .S4_QKV_23(result_QKV_23[59:48]), .S5_QKV_23(result_QKV_23[71:60]), .S6_QKV_23(result_QKV_23[83:72]), .S7_QKV_23(result_QKV_23[95:84]), .S8_QKV_23(result_QKV_23[107:96]), .S9_QKV_23(result_QKV_23[119:108]), .S10_QKV_23(result_QKV_23[131:120]), .S11_QKV_23(result_QKV_23[143:132]), .S12_QKV_23(result_QKV_23[155:144]), .S13_QKV_23(result_QKV_23[167:156]), .S14_QKV_23(result_QKV_23[179:168]), .S15_QKV_23(result_QKV_23[191:180]),
    .S0_QKV_24(result_QKV_24[11:0]), .S1_QKV_24(result_QKV_24[23:12]), .S2_QKV_24(result_QKV_24[35:24]), .S3_QKV_24(result_QKV_24[47:36]), .S4_QKV_24(result_QKV_24[59:48]), .S5_QKV_24(result_QKV_24[71:60]), .S6_QKV_24(result_QKV_24[83:72]), .S7_QKV_24(result_QKV_24[95:84]), .S8_QKV_24(result_QKV_24[107:96]), .S9_QKV_24(result_QKV_24[119:108]), .S10_QKV_24(result_QKV_24[131:120]), .S11_QKV_24(result_QKV_24[143:132]), .S12_QKV_24(result_QKV_24[155:144]), .S13_QKV_24(result_QKV_24[167:156]), .S14_QKV_24(result_QKV_24[179:168]), .S15_QKV_24(result_QKV_24[191:180]),
    .S0_QKV_25(result_QKV_25[11:0]), .S1_QKV_25(result_QKV_25[23:12]), .S2_QKV_25(result_QKV_25[35:24]), .S3_QKV_25(result_QKV_25[47:36]), .S4_QKV_25(result_QKV_25[59:48]), .S5_QKV_25(result_QKV_25[71:60]), .S6_QKV_25(result_QKV_25[83:72]), .S7_QKV_25(result_QKV_25[95:84]), .S8_QKV_25(result_QKV_25[107:96]), .S9_QKV_25(result_QKV_25[119:108]), .S10_QKV_25(result_QKV_25[131:120]), .S11_QKV_25(result_QKV_25[143:132]), .S12_QKV_25(result_QKV_25[155:144]), .S13_QKV_25(result_QKV_25[167:156]), .S14_QKV_25(result_QKV_25[179:168]), .S15_QKV_25(result_QKV_25[191:180]),
    .S0_QKV_26(result_QKV_26[11:0]), .S1_QKV_26(result_QKV_26[23:12]), .S2_QKV_26(result_QKV_26[35:24]), .S3_QKV_26(result_QKV_26[47:36]), .S4_QKV_26(result_QKV_26[59:48]), .S5_QKV_26(result_QKV_26[71:60]), .S6_QKV_26(result_QKV_26[83:72]), .S7_QKV_26(result_QKV_26[95:84]), .S8_QKV_26(result_QKV_26[107:96]), .S9_QKV_26(result_QKV_26[119:108]), .S10_QKV_26(result_QKV_26[131:120]), .S11_QKV_26(result_QKV_26[143:132]), .S12_QKV_26(result_QKV_26[155:144]), .S13_QKV_26(result_QKV_26[167:156]), .S14_QKV_26(result_QKV_26[179:168]), .S15_QKV_26(result_QKV_26[191:180]),
    .S0_QKV_27(result_QKV_27[11:0]), .S1_QKV_27(result_QKV_27[23:12]), .S2_QKV_27(result_QKV_27[35:24]), .S3_QKV_27(result_QKV_27[47:36]), .S4_QKV_27(result_QKV_27[59:48]), .S5_QKV_27(result_QKV_27[71:60]), .S6_QKV_27(result_QKV_27[83:72]), .S7_QKV_27(result_QKV_27[95:84]), .S8_QKV_27(result_QKV_27[107:96]), .S9_QKV_27(result_QKV_27[119:108]), .S10_QKV_27(result_QKV_27[131:120]), .S11_QKV_27(result_QKV_27[143:132]), .S12_QKV_27(result_QKV_27[155:144]), .S13_QKV_27(result_QKV_27[167:156]), .S14_QKV_27(result_QKV_27[179:168]), .S15_QKV_27(result_QKV_27[191:180]),
    .S0_QKV_28(result_QKV_28[11:0]), .S1_QKV_28(result_QKV_28[23:12]), .S2_QKV_28(result_QKV_28[35:24]), .S3_QKV_28(result_QKV_28[47:36]), .S4_QKV_28(result_QKV_28[59:48]), .S5_QKV_28(result_QKV_28[71:60]), .S6_QKV_28(result_QKV_28[83:72]), .S7_QKV_28(result_QKV_28[95:84]), .S8_QKV_28(result_QKV_28[107:96]), .S9_QKV_28(result_QKV_28[119:108]), .S10_QKV_28(result_QKV_28[131:120]), .S11_QKV_28(result_QKV_28[143:132]), .S12_QKV_28(result_QKV_28[155:144]), .S13_QKV_28(result_QKV_28[167:156]), .S14_QKV_28(result_QKV_28[179:168]), .S15_QKV_28(result_QKV_28[191:180]),
    .S0_QKV_29(result_QKV_29[11:0]), .S1_QKV_29(result_QKV_29[23:12]), .S2_QKV_29(result_QKV_29[35:24]), .S3_QKV_29(result_QKV_29[47:36]), .S4_QKV_29(result_QKV_29[59:48]), .S5_QKV_29(result_QKV_29[71:60]), .S6_QKV_29(result_QKV_29[83:72]), .S7_QKV_29(result_QKV_29[95:84]), .S8_QKV_29(result_QKV_29[107:96]), .S9_QKV_29(result_QKV_29[119:108]), .S10_QKV_29(result_QKV_29[131:120]), .S11_QKV_29(result_QKV_29[143:132]), .S12_QKV_29(result_QKV_29[155:144]), .S13_QKV_29(result_QKV_29[167:156]), .S14_QKV_29(result_QKV_29[179:168]), .S15_QKV_29(result_QKV_29[191:180]),
    .S0_QKV_30(result_QKV_30[11:0]), .S1_QKV_30(result_QKV_30[23:12]), .S2_QKV_30(result_QKV_30[35:24]), .S3_QKV_30(result_QKV_30[47:36]), .S4_QKV_30(result_QKV_30[59:48]), .S5_QKV_30(result_QKV_30[71:60]), .S6_QKV_30(result_QKV_30[83:72]), .S7_QKV_30(result_QKV_30[95:84]), .S8_QKV_30(result_QKV_30[107:96]), .S9_QKV_30(result_QKV_30[119:108]), .S10_QKV_30(result_QKV_30[131:120]), .S11_QKV_30(result_QKV_30[143:132]), .S12_QKV_30(result_QKV_30[155:144]), .S13_QKV_30(result_QKV_30[167:156]), .S14_QKV_30(result_QKV_30[179:168]), .S15_QKV_30(result_QKV_30[191:180]),
    .S0_QKV_31(result_QKV_31[11:0]), .S1_QKV_31(result_QKV_31[23:12]), .S2_QKV_31(result_QKV_31[35:24]), .S3_QKV_31(result_QKV_31[47:36]), .S4_QKV_31(result_QKV_31[59:48]), .S5_QKV_31(result_QKV_31[71:60]), .S6_QKV_31(result_QKV_31[83:72]), .S7_QKV_31(result_QKV_31[95:84]), .S8_QKV_31(result_QKV_31[107:96]), .S9_QKV_31(result_QKV_31[119:108]), .S10_QKV_31(result_QKV_31[131:120]), .S11_QKV_31(result_QKV_31[143:132]), .S12_QKV_31(result_QKV_31[155:144]), .S13_QKV_31(result_QKV_31[167:156]), .S14_QKV_31(result_QKV_31[179:168]), .S15_QKV_31(result_QKV_31[191:180]),
    .S0_QKT_0(result_QKT_0[11:0]), .S1_QKT_0(result_QKT_0[23:12]), .S2_QKT_0(result_QKT_0[35:24]), .S3_QKT_0(result_QKT_0[47:36]), .S4_QKT_0(result_QKT_0[59:48]), .S5_QKT_0(result_QKT_0[71:60]), .S6_QKT_0(result_QKT_0[83:72]), .S7_QKT_0(result_QKT_0[95:84]), .S8_QKT_0(result_QKT_0[107:96]), .S9_QKT_0(result_QKT_0[119:108]), .S10_QKT_0(result_QKT_0[131:120]), .S11_QKT_0(result_QKT_0[143:132]), .S12_QKT_0(result_QKT_0[155:144]), .S13_QKT_0(result_QKT_0[167:156]), .S14_QKT_0(result_QKT_0[179:168]), .S15_QKT_0(result_QKT_0[191:180]),
    .S0_QKT_1(result_QKT_1[11:0]), .S1_QKT_1(result_QKT_1[23:12]), .S2_QKT_1(result_QKT_1[35:24]), .S3_QKT_1(result_QKT_1[47:36]), .S4_QKT_1(result_QKT_1[59:48]), .S5_QKT_1(result_QKT_1[71:60]), .S6_QKT_1(result_QKT_1[83:72]), .S7_QKT_1(result_QKT_1[95:84]), .S8_QKT_1(result_QKT_1[107:96]), .S9_QKT_1(result_QKT_1[119:108]), .S10_QKT_1(result_QKT_1[131:120]), .S11_QKT_1(result_QKT_1[143:132]), .S12_QKT_1(result_QKT_1[155:144]), .S13_QKT_1(result_QKT_1[167:156]), .S14_QKT_1(result_QKT_1[179:168]), .S15_QKT_1(result_QKT_1[191:180]),
    .S0_QKT_2(result_QKT_2[11:0]), .S1_QKT_2(result_QKT_2[23:12]), .S2_QKT_2(result_QKT_2[35:24]), .S3_QKT_2(result_QKT_2[47:36]), .S4_QKT_2(result_QKT_2[59:48]), .S5_QKT_2(result_QKT_2[71:60]), .S6_QKT_2(result_QKT_2[83:72]), .S7_QKT_2(result_QKT_2[95:84]), .S8_QKT_2(result_QKT_2[107:96]), .S9_QKT_2(result_QKT_2[119:108]), .S10_QKT_2(result_QKT_2[131:120]), .S11_QKT_2(result_QKT_2[143:132]), .S12_QKT_2(result_QKT_2[155:144]), .S13_QKT_2(result_QKT_2[167:156]), .S14_QKT_2(result_QKT_2[179:168]), .S15_QKT_2(result_QKT_2[191:180]),
    .S0_QKT_3(result_QKT_3[11:0]), .S1_QKT_3(result_QKT_3[23:12]), .S2_QKT_3(result_QKT_3[35:24]), .S3_QKT_3(result_QKT_3[47:36]), .S4_QKT_3(result_QKT_3[59:48]), .S5_QKT_3(result_QKT_3[71:60]), .S6_QKT_3(result_QKT_3[83:72]), .S7_QKT_3(result_QKT_3[95:84]), .S8_QKT_3(result_QKT_3[107:96]), .S9_QKT_3(result_QKT_3[119:108]), .S10_QKT_3(result_QKT_3[131:120]), .S11_QKT_3(result_QKT_3[143:132]), .S12_QKT_3(result_QKT_3[155:144]), .S13_QKT_3(result_QKT_3[167:156]), .S14_QKT_3(result_QKT_3[179:168]), .S15_QKT_3(result_QKT_3[191:180]),


    .WL_QKV_0(WL_QKV_0), .WL_QKV_1(WL_QKV_1), .WL_QKV_2(WL_QKV_2), .WL_QKV_3(WL_QKV_3), .WL_QKV_4(WL_QKV_4), .WL_QKV_5(WL_QKV_5), .WL_QKV_6(WL_QKV_6), .WL_QKV_7(WL_QKV_7), .WL_QKV_8(WL_QKV_8), .WL_QKV_9(WL_QKV_9), .WL_QKV_10(WL_QKV_10), .WL_QKV_11(WL_QKV_11), .WL_QKV_12(WL_QKV_12), .WL_QKV_13(WL_QKV_13), .WL_QKV_14(WL_QKV_14), .WL_QKV_15(WL_QKV_15),
    .WL_QKV_16(WL_QKV_16), .WL_QKV_17(WL_QKV_17), .WL_QKV_18(WL_QKV_18), .WL_QKV_19(WL_QKV_19), .WL_QKV_20(WL_QKV_20), .WL_QKV_21(WL_QKV_21), .WL_QKV_22(WL_QKV_22), .WL_QKV_23(WL_QKV_23), .WL_QKV_24(WL_QKV_24), .WL_QKV_25(WL_QKV_25), .WL_QKV_26(WL_QKV_26), .WL_QKV_27(WL_QKV_27), .WL_QKV_28(WL_QKV_28), .WL_QKV_29(WL_QKV_29), .WL_QKV_30(WL_QKV_30), .WL_QKV_31(WL_QKV_31),
    .WL_QKT_0(WL_QKT_0), .WL_QKT_1(WL_QKT_1), .WL_QKT_2(WL_QKT_2), .WL_QKT_3(WL_QKT_3),

    .wdata_QKV_0(wdata_QKV_0), .wdata_QKV_1(wdata_QKV_1), .wdata_QKV_2(wdata_QKV_2), .wdata_QKV_3(wdata_QKV_3), .wdata_QKV_4(wdata_QKV_4), .wdata_QKV_5(wdata_QKV_5), .wdata_QKV_6(wdata_QKV_6), .wdata_QKV_7(wdata_QKV_7), .wdata_QKV_8(wdata_QKV_8), .wdata_QKV_9(wdata_QKV_9), .wdata_QKV_10(wdata_QKV_10), .wdata_QKV_11(wdata_QKV_11), .wdata_QKV_12(wdata_QKV_12), .wdata_QKV_13(wdata_QKV_13), .wdata_QKV_14(wdata_QKV_14), .wdata_QKV_15(wdata_QKV_15),
    .wdata_QKV_16(wdata_QKV_16), .wdata_QKV_17(wdata_QKV_17), .wdata_QKV_18(wdata_QKV_18), .wdata_QKV_19(wdata_QKV_19), .wdata_QKV_20(wdata_QKV_20), .wdata_QKV_21(wdata_QKV_21), .wdata_QKV_22(wdata_QKV_22), .wdata_QKV_23(wdata_QKV_23), .wdata_QKV_24(wdata_QKV_24), .wdata_QKV_25(wdata_QKV_25), .wdata_QKV_26(wdata_QKV_26), .wdata_QKV_27(wdata_QKV_27), .wdata_QKV_28(wdata_QKV_28), .wdata_QKV_29(wdata_QKV_29), .wdata_QKV_30(wdata_QKV_30), .wdata_QKV_31(wdata_QKV_31),
    .wdata_QKT_0(wdata_QKT_0), .wdata_QKT_1(wdata_QKT_1), .wdata_QKT_2(wdata_QKT_2), .wdata_QKT_3(wdata_QKT_3),

    .ai_QKV_0(ai_QKV_0), .ai_QKV_1(ai_QKV_1), .ai_QKV_2(ai_QKV_2), .ai_QKV_3(ai_QKV_3), .ai_QKV_4(ai_QKV_4), .ai_QKV_5(ai_QKV_5), .ai_QKV_6(ai_QKV_6), .ai_QKV_7(ai_QKV_7), .ai_QKV_8(ai_QKV_8), .ai_QKV_9(ai_QKV_9), .ai_QKV_10(ai_QKV_10), .ai_QKV_11(ai_QKV_11), .ai_QKV_12(ai_QKV_12), .ai_QKV_13(ai_QKV_13), .ai_QKV_14(ai_QKV_14), .ai_QKV_15(ai_QKV_15),
    .ai_QKV_16(ai_QKV_16), .ai_QKV_17(ai_QKV_17), .ai_QKV_18(ai_QKV_18), .ai_QKV_19(ai_QKV_19), .ai_QKV_20(ai_QKV_20), .ai_QKV_21(ai_QKV_21), .ai_QKV_22(ai_QKV_22), .ai_QKV_23(ai_QKV_23), .ai_QKV_24(ai_QKV_24), .ai_QKV_25(ai_QKV_25), .ai_QKV_26(ai_QKV_26), .ai_QKV_27(ai_QKV_27), .ai_QKV_28(ai_QKV_28), .ai_QKV_29(ai_QKV_29), .ai_QKV_30(ai_QKV_30), .ai_QKV_31(ai_QKV_31),
    .ai_QKT_0(ai_QKT_0), .ai_QKT_1(ai_QKT_1), .ai_QKT_2(ai_QKT_2), .ai_QKT_3(ai_QKT_3),

    .RE_QKV__0(RE_QKV__0), .RE_QKV__1(RE_QKV__1), .RE_QKV__2(RE_QKV__2), .RE_QKV__3(RE_QKV__3), .RE_QKV__4(RE_QKV__4), .RE_QKV__5(RE_QKV__5), .RE_QKV__6(RE_QKV__6), .RE_QKV__7(RE_QKV__7), .RE_QKV__8(RE_QKV__8), .RE_QKV__9(RE_QKV__9), .RE_QKV__10(RE_QKV__10), .RE_QKV__11(RE_QKV__11), .RE_QKV__12(RE_QKV__12), .RE_QKV__13(RE_QKV__13), .RE_QKV__14(RE_QKV__14), .RE_QKV__15(RE_QKV__15),
    .RE_QKV__16(RE_QKV__16), .RE_QKV__17(RE_QKV__17), .RE_QKV__18(RE_QKV__18), .RE_QKV__19(RE_QKV__19), .RE_QKV__20(RE_QKV__20), .RE_QKV__21(RE_QKV__21), .RE_QKV__22(RE_QKV__22), .RE_QKV__23(RE_QKV__23), .RE_QKV__24(RE_QKV__24), .RE_QKV__25(RE_QKV__25), .RE_QKV__26(RE_QKV__26), .RE_QKV__27(RE_QKV__27), .RE_QKV__28(RE_QKV__28), .RE_QKV__29(RE_QKV__29), .RE_QKV__30(RE_QKV__30), .RE_QKV__31(RE_QKV__31),
    .RE_QKT__0(RE_QKT__0), .RE_QKT__1(RE_QKT__1), .RE_QKT__2(RE_QKT__2), .RE_QKT__3(RE_QKT__3),

    .PREC_QKV_0(PREC_QKV_0), .PREC_QKV_1(PREC_QKV_1), .PREC_QKV_2(PREC_QKV_2), .PREC_QKV_3(PREC_QKV_3), .PREC_QKV_4(PREC_QKV_4), .PREC_QKV_5(PREC_QKV_5), .PREC_QKV_6(PREC_QKV_6), .PREC_QKV_7(PREC_QKV_7), .PREC_QKV_8(PREC_QKV_8), .PREC_QKV_9(PREC_QKV_9), .PREC_QKV_10(PREC_QKV_10), .PREC_QKV_11(PREC_QKV_11), .PREC_QKV_12(PREC_QKV_12), .PREC_QKV_13(PREC_QKV_13), .PREC_QKV_14(PREC_QKV_14), .PREC_QKV_15(PREC_QKV_15),
    .PREC_QKV_16(PREC_QKV_16), .PREC_QKV_17(PREC_QKV_17), .PREC_QKV_18(PREC_QKV_18), .PREC_QKV_19(PREC_QKV_19), .PREC_QKV_20(PREC_QKV_20), .PREC_QKV_21(PREC_QKV_21), .PREC_QKV_22(PREC_QKV_22), .PREC_QKV_23(PREC_QKV_23), .PREC_QKV_24(PREC_QKV_24), .PREC_QKV_25(PREC_QKV_25), .PREC_QKV_26(PREC_QKV_26), .PREC_QKV_27(PREC_QKV_27), .PREC_QKV_28(PREC_QKV_28), .PREC_QKV_29(PREC_QKV_29), .PREC_QKV_30(PREC_QKV_30), .PREC_QKV_31(PREC_QKV_31),
    .PREC_QKT_0(PREC_QKT_0), .PREC_QKT_1(PREC_QKT_1), .PREC_QKT_2(PREC_QKT_2), .PREC_QKT_3(PREC_QKT_3),

    .PREC_QKV__0(PREC_QKV__0), .PREC_QKV__1(PREC_QKV__1), .PREC_QKV__2(PREC_QKV__2), .PREC_QKV__3(PREC_QKV__3), .PREC_QKV__4(PREC_QKV__4), .PREC_QKV__5(PREC_QKV__5), .PREC_QKV__6(PREC_QKV__6), .PREC_QKV__7(PREC_QKV__7), .PREC_QKV__8(PREC_QKV__8), .PREC_QKV__9(PREC_QKV__9), .PREC_QKV__10(PREC_QKV__10), .PREC_QKV__11(PREC_QKV__11), .PREC_QKV__12(PREC_QKV__12), .PREC_QKV__13(PREC_QKV__13), .PREC_QKV__14(PREC_QKV__14), .PREC_QKV__15(PREC_QKV__15),
    .PREC_QKV__16(PREC_QKV__16), .PREC_QKV__17(PREC_QKV__17), .PREC_QKV__18(PREC_QKV__18), .PREC_QKV__19(PREC_QKV__19), .PREC_QKV__20(PREC_QKV__20), .PREC_QKV__21(PREC_QKV__21), .PREC_QKV__22(PREC_QKV__22), .PREC_QKV__23(PREC_QKV__23), .PREC_QKV__24(PREC_QKV__24), .PREC_QKV__25(PREC_QKV__25), .PREC_QKV__26(PREC_QKV__26), .PREC_QKV__27(PREC_QKV__27), .PREC_QKV__28(PREC_QKV__28), .PREC_QKV__29(PREC_QKV__29), .PREC_QKV__30(PREC_QKV__30), .PREC_QKV__31(PREC_QKV__31),
    .PREC_QKT__0(PREC_QKT__0), .PREC_QKT__1(PREC_QKT__1), .PREC_QKT__2(PREC_QKT__2), .PREC_QKT__3(PREC_QKT__3)
);

`ifdef TARGET_TECH_CELLS_GENERIC_EXCLUDE_TC_SRAM

dimc_macro i_dimc_macro_0(.clk(clk_i),
                          .WL(WL_QKV_0), 
                          .wdata(wdata_QKV_0), 
                          .ai(ai_QKV_0), 
                          .RE_(RE_QKV__0), 
                          .PREC(PREC_QKV_0),
                          .PREC_(PREC_QKV__0),
                          .S0(result_QKV_0[11:0]), 
                          .S1(result_QKV_0[23:12]), 
                          .S2(result_QKV_0[35:24]), 
                          .S3(result_QKV_0[47:36]), 
                          .S4(result_QKV_0[59:48]), 
                          .S5(result_QKV_0[71:60]), 
                          .S6(result_QKV_0[83:72]), 
                          .S7(result_QKV_0[95:84]), 
                          .S8(result_QKV_0[107:96]), 
                          .S9(result_QKV_0[119:108]), 
                          .S10(result_QKV_0[131:120]), 
                          .S11(result_QKV_0[143:132]), 
                          .S12(result_QKV_0[155:144]), 
                          .S13(result_QKV_0[167:156]), 
                          .S14(result_QKV_0[179:168]), 
                          .S15(result_QKV_0[191:180])
                        );

dimc_macro i_dimc_macro_1(.clk(clk_i),
                          .WL(WL_QKV_1), 
                          .wdata(wdata_QKV_1), 
                          .ai(ai_QKV_1), 
                          .RE_(RE_QKV__1), 
                          .PREC(PREC_QKV_1),
                          .PREC_(PREC_QKV__1),
                          .S0(result_QKV_1[11:0]), 
                          .S1(result_QKV_1[23:12]), 
                          .S2(result_QKV_1[35:24]), 
                          .S3(result_QKV_1[47:36]), 
                          .S4(result_QKV_1[59:48]), 
                          .S5(result_QKV_1[71:60]), 
                          .S6(result_QKV_1[83:72]), 
                          .S7(result_QKV_1[95:84]), 
                          .S8(result_QKV_1[107:96]), 
                          .S9(result_QKV_1[119:108]), 
                          .S10(result_QKV_1[131:120]), 
                          .S11(result_QKV_1[143:132]), 
                          .S12(result_QKV_1[155:144]), 
                          .S13(result_QKV_1[167:156]), 
                          .S14(result_QKV_1[179:168]), 
                          .S15(result_QKV_1[191:180])
                        );

dimc_macro i_dimc_macro_2(.clk(clk_i),
                          .WL(WL_QKV_2), 
                          .wdata(wdata_QKV_2), 
                          .ai(ai_QKV_2), 
                          .RE_(RE_QKV__2), 
                          .PREC(PREC_QKV_2),
                          .PREC_(PREC_QKV__2),
                          .S0(result_QKV_2[11:0]), 
                          .S1(result_QKV_2[23:12]), 
                          .S2(result_QKV_2[35:24]), 
                          .S3(result_QKV_2[47:36]), 
                          .S4(result_QKV_2[59:48]), 
                          .S5(result_QKV_2[71:60]), 
                          .S6(result_QKV_2[83:72]), 
                          .S7(result_QKV_2[95:84]), 
                          .S8(result_QKV_2[107:96]), 
                          .S9(result_QKV_2[119:108]), 
                          .S10(result_QKV_2[131:120]), 
                          .S11(result_QKV_2[143:132]), 
                          .S12(result_QKV_2[155:144]), 
                          .S13(result_QKV_2[167:156]), 
                          .S14(result_QKV_2[179:168]), 
                          .S15(result_QKV_2[191:180])
                        );

dimc_macro i_dimc_macro_3(.clk(clk_i),
                          .WL(WL_QKV_3), 
                          .wdata(wdata_QKV_3), 
                          .ai(ai_QKV_3), 
                          .RE_(RE_QKV__3), 
                          .PREC(PREC_QKV_3),
                          .PREC_(PREC_QKV__3),
                          .S0(result_QKV_3[11:0]),
                          .S1(result_QKV_3[23:12]),
                          .S2(result_QKV_3[35:24]),
                          .S3(result_QKV_3[47:36]),
                          .S4(result_QKV_3[59:48]),
                          .S5(result_QKV_3[71:60]),
                          .S6(result_QKV_3[83:72]),
                          .S7(result_QKV_3[95:84]),
                          .S8(result_QKV_3[107:96]),
                          .S9(result_QKV_3[119:108]),
                          .S10(result_QKV_3[131:120]),
                          .S11(result_QKV_3[143:132]),
                          .S12(result_QKV_3[155:144]),
                          .S13(result_QKV_3[167:156]),
                          .S14(result_QKV_3[179:168]),
                          .S15(result_QKV_3[191:180])
                        );

dimc_macro i_dimc_macro_4(.clk(clk_i),
                          .WL(WL_QKV_4), 
                          .wdata(wdata_QKV_4), 
                          .ai(ai_QKV_4), 
                          .RE_(RE_QKV__4), 
                          .PREC(PREC_QKV_4),
                          .PREC_(PREC_QKV__4),
                          .S0(result_QKV_4[11:0]), 
                          .S1(result_QKV_4[23:12]), 
                          .S2(result_QKV_4[35:24]), 
                          .S3(result_QKV_4[47:36]), 
                          .S4(result_QKV_4[59:48]), 
                          .S5(result_QKV_4[71:60]), 
                          .S6(result_QKV_4[83:72]), 
                          .S7(result_QKV_4[95:84]), 
                          .S8(result_QKV_4[107:96]), 
                          .S9(result_QKV_4[119:108]), 
                          .S10(result_QKV_4[131:120]), 
                          .S11(result_QKV_4[143:132]), 
                          .S12(result_QKV_4[155:144]), 
                          .S13(result_QKV_4[167:156]), 
                          .S14(result_QKV_4[179:168]), 
                          .S15(result_QKV_4[191:180])
                        );

dimc_macro i_dimc_macro_5(.clk(clk_i),
                          .WL(WL_QKV_5), 
                          .wdata(wdata_QKV_5), 
                          .ai(ai_QKV_5), 
                          .RE_(RE_QKV__5), 
                          .PREC(PREC_QKV_5),
                          .PREC_(PREC_QKV__5),
                          .S0(result_QKV_5[11:0]), 
                          .S1(result_QKV_5[23:12]), 
                          .S2(result_QKV_5[35:24]), 
                          .S3(result_QKV_5[47:36]), 
                          .S4(result_QKV_5[59:48]), 
                          .S5(result_QKV_5[71:60]), 
                          .S6(result_QKV_5[83:72]), 
                          .S7(result_QKV_5[95:84]), 
                          .S8(result_QKV_5[107:96]), 
                          .S9(result_QKV_5[119:108]), 
                          .S10(result_QKV_5[131:120]), 
                          .S11(result_QKV_5[143:132]), 
                          .S12(result_QKV_5[155:144]), 
                          .S13(result_QKV_5[167:156]), 
                          .S14(result_QKV_5[179:168]), 
                          .S15(result_QKV_5[191:180])
                        );

dimc_macro i_dimc_macro_6(.clk(clk_i),
                          .WL(WL_QKV_6), 
                          .wdata(wdata_QKV_6), 
                          .ai(ai_QKV_6), 
                          .RE_(RE_QKV__6), 
                          .PREC(PREC_QKV_6),
                          .PREC_(PREC_QKV__6),
                          .S0(result_QKV_6[11:0]), 
                          .S1(result_QKV_6[23:12]), 
                          .S2(result_QKV_6[35:24]), 
                          .S3(result_QKV_6[47:36]), 
                          .S4(result_QKV_6[59:48]), 
                          .S5(result_QKV_6[71:60]), 
                          .S6(result_QKV_6[83:72]), 
                          .S7(result_QKV_6[95:84]), 
                          .S8(result_QKV_6[107:96]), 
                          .S9(result_QKV_6[119:108]), 
                          .S10(result_QKV_6[131:120]), 
                          .S11(result_QKV_6[143:132]), 
                          .S12(result_QKV_6[155:144]), 
                          .S13(result_QKV_6[167:156]), 
                          .S14(result_QKV_6[179:168]), 
                          .S15(result_QKV_6[191:180])
                        );

dimc_macro i_dimc_macro_7(.clk(clk_i),
                          .WL(WL_QKV_7), 
                          .wdata(wdata_QKV_7), 
                          .ai(ai_QKV_7), 
                          .RE_(RE_QKV__7), 
                          .PREC(PREC_QKV_7),
                          .PREC_(PREC_QKV__7),
                          .S0(result_QKV_7[11:0]), 
                          .S1(result_QKV_7[23:12]), 
                          .S2(result_QKV_7[35:24]), 
                          .S3(result_QKV_7[47:36]), 
                          .S4(result_QKV_7[59:48]), 
                          .S5(result_QKV_7[71:60]), 
                          .S6(result_QKV_7[83:72]), 
                          .S7(result_QKV_7[95:84]), 
                          .S8(result_QKV_7[107:96]), 
                          .S9(result_QKV_7[119:108]), 
                          .S10(result_QKV_7[131:120]), 
                          .S11(result_QKV_7[143:132]), 
                          .S12(result_QKV_7[155:144]), 
                          .S13(result_QKV_7[167:156]), 
                          .S14(result_QKV_7[179:168]), 
                          .S15(result_QKV_7[191:180])
                        );

dimc_macro i_dimc_macro_8(.clk(clk_i),
                          .WL(WL_QKV_8), 
                          .wdata(wdata_QKV_8), 
                          .ai(ai_QKV_8), 
                          .RE_(RE_QKV__8), 
                          .PREC(PREC_QKV_8),
                          .PREC_(PREC_QKV__8),
                          .S0(result_QKV_8[11:0]), 
                          .S1(result_QKV_8[23:12]), 
                          .S2(result_QKV_8[35:24]), 
                          .S3(result_QKV_8[47:36]), 
                          .S4(result_QKV_8[59:48]), 
                          .S5(result_QKV_8[71:60]), 
                          .S6(result_QKV_8[83:72]), 
                          .S7(result_QKV_8[95:84]), 
                          .S8(result_QKV_8[107:96]), 
                          .S9(result_QKV_8[119:108]), 
                          .S10(result_QKV_8[131:120]), 
                          .S11(result_QKV_8[143:132]), 
                          .S12(result_QKV_8[155:144]), 
                          .S13(result_QKV_8[167:156]), 
                          .S14(result_QKV_8[179:168]), 
                          .S15(result_QKV_8[191:180])
                        );

dimc_macro i_dimc_macro_9(.clk(clk_i),
                          .WL(WL_QKV_9), 
                          .wdata(wdata_QKV_9), 
                          .ai(ai_QKV_9), 
                          .RE_(RE_QKV__9), 
                          .PREC(PREC_QKV_9),
                          .PREC_(PREC_QKV__9),
                          .S0(result_QKV_9[11:0]), 
                          .S1(result_QKV_9[23:12]), 
                          .S2(result_QKV_9[35:24]), 
                          .S3(result_QKV_9[47:36]), 
                          .S4(result_QKV_9[59:48]), 
                          .S5(result_QKV_9[71:60]), 
                          .S6(result_QKV_9[83:72]), 
                          .S7(result_QKV_9[95:84]), 
                          .S8(result_QKV_9[107:96]), 
                          .S9(result_QKV_9[119:108]), 
                          .S10(result_QKV_9[131:120]), 
                          .S11(result_QKV_9[143:132]), 
                          .S12(result_QKV_9[155:144]), 
                          .S13(result_QKV_9[167:156]), 
                          .S14(result_QKV_9[179:168]), 
                          .S15(result_QKV_9[191:180])
                        );

dimc_macro i_dimc_macro_10(.clk(clk_i),
                          .WL(WL_QKV_10), 
                          .wdata(wdata_QKV_10), 
                          .ai(ai_QKV_10), 
                          .RE_(RE_QKV__10), 
                          .PREC(PREC_QKV_10),
                          .PREC_(PREC_QKV__10),
                          .S0(result_QKV_10[11:0]), 
                          .S1(result_QKV_10[23:12]), 
                          .S2(result_QKV_10[35:24]), 
                          .S3(result_QKV_10[47:36]), 
                          .S4(result_QKV_10[59:48]), 
                          .S5(result_QKV_10[71:60]), 
                          .S6(result_QKV_10[83:72]), 
                          .S7(result_QKV_10[95:84]), 
                          .S8(result_QKV_10[107:96]), 
                          .S9(result_QKV_10[119:108]), 
                          .S10(result_QKV_10[131:120]), 
                          .S11(result_QKV_10[143:132]), 
                          .S12(result_QKV_10[155:144]), 
                          .S13(result_QKV_10[167:156]), 
                          .S14(result_QKV_10[179:168]), 
                          .S15(result_QKV_10[191:180])
                        );

dimc_macro i_dimc_macro_11(.clk(clk_i),
                          .WL(WL_QKV_11), 
                          .wdata(wdata_QKV_11), 
                          .ai(ai_QKV_11), 
                          .RE_(RE_QKV__11), 
                          .PREC(PREC_QKV_11),
                          .PREC_(PREC_QKV__11),
                          .S0(result_QKV_11[11:0]), 
                          .S1(result_QKV_11[23:12]), 
                          .S2(result_QKV_11[35:24]), 
                          .S3(result_QKV_11[47:36]), 
                          .S4(result_QKV_11[59:48]), 
                          .S5(result_QKV_11[71:60]), 
                          .S6(result_QKV_11[83:72]), 
                          .S7(result_QKV_11[95:84]), 
                          .S8(result_QKV_11[107:96]), 
                          .S9(result_QKV_11[119:108]), 
                          .S10(result_QKV_11[131:120]), 
                          .S11(result_QKV_11[143:132]), 
                          .S12(result_QKV_11[155:144]), 
                          .S13(result_QKV_11[167:156]), 
                          .S14(result_QKV_11[179:168]), 
                          .S15(result_QKV_11[191:180])
                        );

dimc_macro i_dimc_macro_12(.clk(clk_i),
                          .WL(WL_QKV_12), 
                          .wdata(wdata_QKV_12), 
                          .ai(ai_QKV_12), 
                          .RE_(RE_QKV__12), 
                          .PREC(PREC_QKV_12),
                          .PREC_(PREC_QKV__12),
                          .S0(result_QKV_12[11:0]), 
                          .S1(result_QKV_12[23:12]), 
                          .S2(result_QKV_12[35:24]), 
                          .S3(result_QKV_12[47:36]), 
                          .S4(result_QKV_12[59:48]), 
                          .S5(result_QKV_12[71:60]), 
                          .S6(result_QKV_12[83:72]), 
                          .S7(result_QKV_12[95:84]), 
                          .S8(result_QKV_12[107:96]), 
                          .S9(result_QKV_12[119:108]), 
                          .S10(result_QKV_12[131:120]), 
                          .S11(result_QKV_12[143:132]), 
                          .S12(result_QKV_12[155:144]), 
                          .S13(result_QKV_12[167:156]), 
                          .S14(result_QKV_12[179:168]), 
                          .S15(result_QKV_12[191:180])
                        );

dimc_macro i_dimc_macro_13(.clk(clk_i),
                          .WL(WL_QKV_13), 
                          .wdata(wdata_QKV_13), 
                          .ai(ai_QKV_13), 
                          .RE_(RE_QKV__13), 
                          .PREC(PREC_QKV_13),
                          .PREC_(PREC_QKV__13),
                          .S0(result_QKV_13[11:0]), 
                          .S1(result_QKV_13[23:12]), 
                          .S2(result_QKV_13[35:24]), 
                          .S3(result_QKV_13[47:36]), 
                          .S4(result_QKV_13[59:48]), 
                          .S5(result_QKV_13[71:60]), 
                          .S6(result_QKV_13[83:72]), 
                          .S7(result_QKV_13[95:84]), 
                          .S8(result_QKV_13[107:96]), 
                          .S9(result_QKV_13[119:108]), 
                          .S10(result_QKV_13[131:120]), 
                          .S11(result_QKV_13[143:132]), 
                          .S12(result_QKV_13[155:144]), 
                          .S13(result_QKV_13[167:156]), 
                          .S14(result_QKV_13[179:168]), 
                          .S15(result_QKV_13[191:180])
                        );

dimc_macro i_dimc_macro_14(.clk(clk_i),
                          .WL(WL_QKV_14), 
                          .wdata(wdata_QKV_14), 
                          .ai(ai_QKV_14), 
                          .RE_(RE_QKV__14), 
                          .PREC(PREC_QKV_14),
                          .PREC_(PREC_QKV__14),
                          .S0(result_QKV_14[11:0]), 
                          .S1(result_QKV_14[23:12]), 
                          .S2(result_QKV_14[35:24]), 
                          .S3(result_QKV_14[47:36]), 
                          .S4(result_QKV_14[59:48]), 
                          .S5(result_QKV_14[71:60]), 
                          .S6(result_QKV_14[83:72]), 
                          .S7(result_QKV_14[95:84]), 
                          .S8(result_QKV_14[107:96]), 
                          .S9(result_QKV_14[119:108]), 
                          .S10(result_QKV_14[131:120]), 
                          .S11(result_QKV_14[143:132]), 
                          .S12(result_QKV_14[155:144]), 
                          .S13(result_QKV_14[167:156]), 
                          .S14(result_QKV_14[179:168]), 
                          .S15(result_QKV_14[191:180])
                        );

dimc_macro i_dimc_macro_15(.clk(clk_i),
                          .WL(WL_QKV_15), 
                          .wdata(wdata_QKV_15), 
                          .ai(ai_QKV_15), 
                          .RE_(RE_QKV__15), 
                          .PREC(PREC_QKV_15),
                          .PREC_(PREC_QKV__15),
                          .S0(result_QKV_15[11:0]), 
                          .S1(result_QKV_15[23:12]), 
                          .S2(result_QKV_15[35:24]), 
                          .S3(result_QKV_15[47:36]), 
                          .S4(result_QKV_15[59:48]), 
                          .S5(result_QKV_15[71:60]), 
                          .S6(result_QKV_15[83:72]), 
                          .S7(result_QKV_15[95:84]), 
                          .S8(result_QKV_15[107:96]), 
                          .S9(result_QKV_15[119:108]), 
                          .S10(result_QKV_15[131:120]), 
                          .S11(result_QKV_15[143:132]), 
                          .S12(result_QKV_15[155:144]), 
                          .S13(result_QKV_15[167:156]), 
                          .S14(result_QKV_15[179:168]), 
                          .S15(result_QKV_15[191:180])
                        );

dimc_macro i_dimc_macro_16(.clk(clk_i),
                          .WL(WL_QKV_16), 
                          .wdata(wdata_QKV_16), 
                          .ai(ai_QKV_16), 
                          .RE_(RE_QKV__16), 
                          .PREC(PREC_QKV_16),
                          .PREC_(PREC_QKV__16),
                          .S0(result_QKV_16[11:0]), 
                          .S1(result_QKV_16[23:12]), 
                          .S2(result_QKV_16[35:24]), 
                          .S3(result_QKV_16[47:36]), 
                          .S4(result_QKV_16[59:48]), 
                          .S5(result_QKV_16[71:60]), 
                          .S6(result_QKV_16[83:72]), 
                          .S7(result_QKV_16[95:84]), 
                          .S8(result_QKV_16[107:96]), 
                          .S9(result_QKV_16[119:108]), 
                          .S10(result_QKV_16[131:120]), 
                          .S11(result_QKV_16[143:132]), 
                          .S12(result_QKV_16[155:144]), 
                          .S13(result_QKV_16[167:156]), 
                          .S14(result_QKV_16[179:168]), 
                          .S15(result_QKV_16[191:180])
                        );

dimc_macro i_dimc_macro_17(.clk(clk_i),
                          .WL(WL_QKV_17), 
                          .wdata(wdata_QKV_17), 
                          .ai(ai_QKV_17), 
                          .RE_(RE_QKV__17), 
                          .PREC(PREC_QKV_17),
                          .PREC_(PREC_QKV__17),
                          .S0(result_QKV_17[11:0]), 
                          .S1(result_QKV_17[23:12]), 
                          .S2(result_QKV_17[35:24]), 
                          .S3(result_QKV_17[47:36]), 
                          .S4(result_QKV_17[59:48]), 
                          .S5(result_QKV_17[71:60]), 
                          .S6(result_QKV_17[83:72]), 
                          .S7(result_QKV_17[95:84]), 
                          .S8(result_QKV_17[107:96]), 
                          .S9(result_QKV_17[119:108]), 
                          .S10(result_QKV_17[131:120]), 
                          .S11(result_QKV_17[143:132]), 
                          .S12(result_QKV_17[155:144]), 
                          .S13(result_QKV_17[167:156]), 
                          .S14(result_QKV_17[179:168]), 
                          .S15(result_QKV_17[191:180])
                        );

dimc_macro i_dimc_macro_18(.clk(clk_i),
                          .WL(WL_QKV_18), 
                          .wdata(wdata_QKV_18), 
                          .ai(ai_QKV_18), 
                          .RE_(RE_QKV__18), 
                          .PREC(PREC_QKV_18),
                          .PREC_(PREC_QKV__18),
                          .S0(result_QKV_18[11:0]), 
                          .S1(result_QKV_18[23:12]), 
                          .S2(result_QKV_18[35:24]), 
                          .S3(result_QKV_18[47:36]), 
                          .S4(result_QKV_18[59:48]), 
                          .S5(result_QKV_18[71:60]), 
                          .S6(result_QKV_18[83:72]), 
                          .S7(result_QKV_18[95:84]), 
                          .S8(result_QKV_18[107:96]), 
                          .S9(result_QKV_18[119:108]), 
                          .S10(result_QKV_18[131:120]), 
                          .S11(result_QKV_18[143:132]), 
                          .S12(result_QKV_18[155:144]), 
                          .S13(result_QKV_18[167:156]), 
                          .S14(result_QKV_18[179:168]), 
                          .S15(result_QKV_18[191:180])
                        );

dimc_macro i_dimc_macro_19(.clk(clk_i),
                          .WL(WL_QKV_19), 
                          .wdata(wdata_QKV_19), 
                          .ai(ai_QKV_19), 
                          .RE_(RE_QKV__19), 
                          .PREC(PREC_QKV_19),
                          .PREC_(PREC_QKV__19),
                          .S0(result_QKV_19[11:0]), 
                          .S1(result_QKV_19[23:12]), 
                          .S2(result_QKV_19[35:24]), 
                          .S3(result_QKV_19[47:36]), 
                          .S4(result_QKV_19[59:48]), 
                          .S5(result_QKV_19[71:60]), 
                          .S6(result_QKV_19[83:72]), 
                          .S7(result_QKV_19[95:84]), 
                          .S8(result_QKV_19[107:96]), 
                          .S9(result_QKV_19[119:108]), 
                          .S10(result_QKV_19[131:120]), 
                          .S11(result_QKV_19[143:132]), 
                          .S12(result_QKV_19[155:144]), 
                          .S13(result_QKV_19[167:156]), 
                          .S14(result_QKV_19[179:168]), 
                          .S15(result_QKV_19[191:180])
                        );

dimc_macro i_dimc_macro_20(.clk(clk_i),
                          .WL(WL_QKV_20), 
                          .wdata(wdata_QKV_20), 
                          .ai(ai_QKV_20), 
                          .RE_(RE_QKV__20), 
                          .PREC(PREC_QKV_20),
                          .PREC_(PREC_QKV__20),
                          .S0(result_QKV_20[11:0]), 
                          .S1(result_QKV_20[23:12]), 
                          .S2(result_QKV_20[35:24]), 
                          .S3(result_QKV_20[47:36]), 
                          .S4(result_QKV_20[59:48]), 
                          .S5(result_QKV_20[71:60]), 
                          .S6(result_QKV_20[83:72]), 
                          .S7(result_QKV_20[95:84]), 
                          .S8(result_QKV_20[107:96]), 
                          .S9(result_QKV_20[119:108]), 
                          .S10(result_QKV_20[131:120]), 
                          .S11(result_QKV_20[143:132]), 
                          .S12(result_QKV_20[155:144]), 
                          .S13(result_QKV_20[167:156]), 
                          .S14(result_QKV_20[179:168]), 
                          .S15(result_QKV_20[191:180])
                        );

dimc_macro i_dimc_macro_21(.clk(clk_i),
                          .WL(WL_QKV_21), 
                          .wdata(wdata_QKV_21), 
                          .ai(ai_QKV_21), 
                          .RE_(RE_QKV__21), 
                          .PREC(PREC_QKV_21),
                          .PREC_(PREC_QKV__21),
                          .S0(result_QKV_21[11:0]), 
                          .S1(result_QKV_21[23:12]), 
                          .S2(result_QKV_21[35:24]), 
                          .S3(result_QKV_21[47:36]), 
                          .S4(result_QKV_21[59:48]), 
                          .S5(result_QKV_21[71:60]), 
                          .S6(result_QKV_21[83:72]), 
                          .S7(result_QKV_21[95:84]), 
                          .S8(result_QKV_21[107:96]), 
                          .S9(result_QKV_21[119:108]), 
                          .S10(result_QKV_21[131:120]), 
                          .S11(result_QKV_21[143:132]), 
                          .S12(result_QKV_21[155:144]), 
                          .S13(result_QKV_21[167:156]), 
                          .S14(result_QKV_21[179:168]), 
                          .S15(result_QKV_21[191:180])
                        );

dimc_macro i_dimc_macro_22(.clk(clk_i),
                          .WL(WL_QKV_22), 
                          .wdata(wdata_QKV_22), 
                          .ai(ai_QKV_22), 
                          .RE_(RE_QKV__22), 
                          .PREC(PREC_QKV_22),
                          .PREC_(PREC_QKV__22),
                          .S0(result_QKV_22[11:0]), 
                          .S1(result_QKV_22[23:12]), 
                          .S2(result_QKV_22[35:24]), 
                          .S3(result_QKV_22[47:36]), 
                          .S4(result_QKV_22[59:48]), 
                          .S5(result_QKV_22[71:60]), 
                          .S6(result_QKV_22[83:72]), 
                          .S7(result_QKV_22[95:84]), 
                          .S8(result_QKV_22[107:96]), 
                          .S9(result_QKV_22[119:108]), 
                          .S10(result_QKV_22[131:120]), 
                          .S11(result_QKV_22[143:132]), 
                          .S12(result_QKV_22[155:144]), 
                          .S13(result_QKV_22[167:156]), 
                          .S14(result_QKV_22[179:168]), 
                          .S15(result_QKV_22[191:180])
                        );

dimc_macro i_dimc_macro_23(.clk(clk_i),
                          .WL(WL_QKV_23), 
                          .wdata(wdata_QKV_23), 
                          .ai(ai_QKV_23), 
                          .RE_(RE_QKV__23), 
                          .PREC(PREC_QKV_23),
                          .PREC_(PREC_QKV__23),
                          .S0(result_QKV_23[11:0]), 
                          .S1(result_QKV_23[23:12]), 
                          .S2(result_QKV_23[35:24]), 
                          .S3(result_QKV_23[47:36]), 
                          .S4(result_QKV_23[59:48]), 
                          .S5(result_QKV_23[71:60]), 
                          .S6(result_QKV_23[83:72]), 
                          .S7(result_QKV_23[95:84]), 
                          .S8(result_QKV_23[107:96]), 
                          .S9(result_QKV_23[119:108]), 
                          .S10(result_QKV_23[131:120]), 
                          .S11(result_QKV_23[143:132]), 
                          .S12(result_QKV_23[155:144]), 
                          .S13(result_QKV_23[167:156]), 
                          .S14(result_QKV_23[179:168]), 
                          .S15(result_QKV_23[191:180])
                        );

dimc_macro i_dimc_macro_24(.clk(clk_i),
                          .WL(WL_QKV_24), 
                          .wdata(wdata_QKV_24), 
                          .ai(ai_QKV_24), 
                          .RE_(RE_QKV__24), 
                          .PREC(PREC_QKV_24),
                          .PREC_(PREC_QKV__24),
                          .S0(result_QKV_24[11:0]), 
                          .S1(result_QKV_24[23:12]), 
                          .S2(result_QKV_24[35:24]), 
                          .S3(result_QKV_24[47:36]), 
                          .S4(result_QKV_24[59:48]), 
                          .S5(result_QKV_24[71:60]), 
                          .S6(result_QKV_24[83:72]), 
                          .S7(result_QKV_24[95:84]), 
                          .S8(result_QKV_24[107:96]), 
                          .S9(result_QKV_24[119:108]), 
                          .S10(result_QKV_24[131:120]), 
                          .S11(result_QKV_24[143:132]), 
                          .S12(result_QKV_24[155:144]), 
                          .S13(result_QKV_24[167:156]), 
                          .S14(result_QKV_24[179:168]), 
                          .S15(result_QKV_24[191:180])
                        );

dimc_macro i_dimc_macro_25(.clk(clk_i),
                          .WL(WL_QKV_25), 
                          .wdata(wdata_QKV_25), 
                          .ai(ai_QKV_25), 
                          .RE_(RE_QKV__25), 
                          .PREC(PREC_QKV_25),
                          .PREC_(PREC_QKV__25),
                          .S0(result_QKV_25[11:0]), 
                          .S1(result_QKV_25[23:12]), 
                          .S2(result_QKV_25[35:24]), 
                          .S3(result_QKV_25[47:36]), 
                          .S4(result_QKV_25[59:48]), 
                          .S5(result_QKV_25[71:60]), 
                          .S6(result_QKV_25[83:72]), 
                          .S7(result_QKV_25[95:84]), 
                          .S8(result_QKV_25[107:96]), 
                          .S9(result_QKV_25[119:108]), 
                          .S10(result_QKV_25[131:120]), 
                          .S11(result_QKV_25[143:132]), 
                          .S12(result_QKV_25[155:144]), 
                          .S13(result_QKV_25[167:156]), 
                          .S14(result_QKV_25[179:168]), 
                          .S15(result_QKV_25[191:180])
                        );

dimc_macro i_dimc_macro_26(.clk(clk_i),
                          .WL(WL_QKV_26), 
                          .wdata(wdata_QKV_26), 
                          .ai(ai_QKV_26), 
                          .RE_(RE_QKV__26), 
                          .PREC(PREC_QKV_26),
                          .PREC_(PREC_QKV__26),
                          .S0(result_QKV_26[11:0]), 
                          .S1(result_QKV_26[23:12]), 
                          .S2(result_QKV_26[35:24]), 
                          .S3(result_QKV_26[47:36]), 
                          .S4(result_QKV_26[59:48]), 
                          .S5(result_QKV_26[71:60]), 
                          .S6(result_QKV_26[83:72]), 
                          .S7(result_QKV_26[95:84]), 
                          .S8(result_QKV_26[107:96]), 
                          .S9(result_QKV_26[119:108]), 
                          .S10(result_QKV_26[131:120]), 
                          .S11(result_QKV_26[143:132]), 
                          .S12(result_QKV_26[155:144]), 
                          .S13(result_QKV_26[167:156]), 
                          .S14(result_QKV_26[179:168]), 
                          .S15(result_QKV_26[191:180])
                        );

dimc_macro i_dimc_macro_27(.clk(clk_i),
                          .WL(WL_QKV_27), 
                          .wdata(wdata_QKV_27), 
                          .ai(ai_QKV_27), 
                          .RE_(RE_QKV__27), 
                          .PREC(PREC_QKV_27),
                          .PREC_(PREC_QKV__27),
                          .S0(result_QKV_27[11:0]), 
                          .S1(result_QKV_27[23:12]), 
                          .S2(result_QKV_27[35:24]), 
                          .S3(result_QKV_27[47:36]), 
                          .S4(result_QKV_27[59:48]), 
                          .S5(result_QKV_27[71:60]), 
                          .S6(result_QKV_27[83:72]), 
                          .S7(result_QKV_27[95:84]), 
                          .S8(result_QKV_27[107:96]), 
                          .S9(result_QKV_27[119:108]), 
                          .S10(result_QKV_27[131:120]), 
                          .S11(result_QKV_27[143:132]), 
                          .S12(result_QKV_27[155:144]), 
                          .S13(result_QKV_27[167:156]), 
                          .S14(result_QKV_27[179:168]), 
                          .S15(result_QKV_27[191:180])
                        );

dimc_macro i_dimc_macro_28(.clk(clk_i),
                          .WL(WL_QKV_28), 
                          .wdata(wdata_QKV_28), 
                          .ai(ai_QKV_28), 
                          .RE_(RE_QKV__28), 
                          .PREC(PREC_QKV_28),
                          .PREC_(PREC_QKV__28),
                          .S0(result_QKV_28[11:0]), 
                          .S1(result_QKV_28[23:12]), 
                          .S2(result_QKV_28[35:24]), 
                          .S3(result_QKV_28[47:36]), 
                          .S4(result_QKV_28[59:48]), 
                          .S5(result_QKV_28[71:60]), 
                          .S6(result_QKV_28[83:72]), 
                          .S7(result_QKV_28[95:84]), 
                          .S8(result_QKV_28[107:96]), 
                          .S9(result_QKV_28[119:108]), 
                          .S10(result_QKV_28[131:120]), 
                          .S11(result_QKV_28[143:132]), 
                          .S12(result_QKV_28[155:144]), 
                          .S13(result_QKV_28[167:156]), 
                          .S14(result_QKV_28[179:168]), 
                          .S15(result_QKV_28[191:180])
                        );

dimc_macro i_dimc_macro_29(.clk(clk_i),
                          .WL(WL_QKV_29), 
                          .wdata(wdata_QKV_29), 
                          .ai(ai_QKV_29), 
                          .RE_(RE_QKV__29), 
                          .PREC(PREC_QKV_29),
                          .PREC_(PREC_QKV__29),
                          .S0(result_QKV_29[11:0]), 
                          .S1(result_QKV_29[23:12]), 
                          .S2(result_QKV_29[35:24]), 
                          .S3(result_QKV_29[47:36]), 
                          .S4(result_QKV_29[59:48]), 
                          .S5(result_QKV_29[71:60]), 
                          .S6(result_QKV_29[83:72]), 
                          .S7(result_QKV_29[95:84]), 
                          .S8(result_QKV_29[107:96]), 
                          .S9(result_QKV_29[119:108]), 
                          .S10(result_QKV_29[131:120]), 
                          .S11(result_QKV_29[143:132]), 
                          .S12(result_QKV_29[155:144]), 
                          .S13(result_QKV_29[167:156]), 
                          .S14(result_QKV_29[179:168]), 
                          .S15(result_QKV_29[191:180])
                        );

dimc_macro i_dimc_macro_30(.clk(clk_i),
                          .WL(WL_QKV_30), 
                          .wdata(wdata_QKV_30), 
                          .ai(ai_QKV_30), 
                          .RE_(RE_QKV__30), 
                          .PREC(PREC_QKV_30),
                          .PREC_(PREC_QKV__30),
                          .S0(result_QKV_30[11:0]), 
                          .S1(result_QKV_30[23:12]), 
                          .S2(result_QKV_30[35:24]), 
                          .S3(result_QKV_30[47:36]), 
                          .S4(result_QKV_30[59:48]), 
                          .S5(result_QKV_30[71:60]), 
                          .S6(result_QKV_30[83:72]), 
                          .S7(result_QKV_30[95:84]), 
                          .S8(result_QKV_30[107:96]), 
                          .S9(result_QKV_30[119:108]), 
                          .S10(result_QKV_30[131:120]), 
                          .S11(result_QKV_30[143:132]), 
                          .S12(result_QKV_30[155:144]), 
                          .S13(result_QKV_30[167:156]), 
                          .S14(result_QKV_30[179:168]), 
                          .S15(result_QKV_30[191:180])
                        );

dimc_macro i_dimc_macro_31(.clk(clk_i),
                          .WL(WL_QKV_31), 
                          .wdata(wdata_QKV_31), 
                          .ai(ai_QKV_31), 
                          .RE_(RE_QKV__31), 
                          .PREC(PREC_QKV_31),
                          .PREC_(PREC_QKV__31),
                          .S0(result_QKV_31[11:0]), 
                          .S1(result_QKV_31[23:12]), 
                          .S2(result_QKV_31[35:24]), 
                          .S3(result_QKV_31[47:36]), 
                          .S4(result_QKV_31[59:48]), 
                          .S5(result_QKV_31[71:60]), 
                          .S6(result_QKV_31[83:72]), 
                          .S7(result_QKV_31[95:84]), 
                          .S8(result_QKV_31[107:96]), 
                          .S9(result_QKV_31[119:108]), 
                          .S10(result_QKV_31[131:120]), 
                          .S11(result_QKV_31[143:132]), 
                          .S12(result_QKV_31[155:144]), 
                          .S13(result_QKV_31[167:156]), 
                          .S14(result_QKV_31[179:168]), 
                          .S15(result_QKV_31[191:180])
                        );

dimc_macro i_dimc_macro_32(.clk(clk_i),
                          .WL(WL_QKT_0), 
                          .wdata(wdata_QKT_0), 
                          .ai(ai_QKT_0), 
                          .RE_(RE_QKT__0), 
                          .PREC(PREC_QKT_0),
                          .PREC_(PREC_QKT__0),
                          .S0(result_QKT_0[11:0]), 
                          .S1(result_QKT_0[23:12]), 
                          .S2(result_QKT_0[35:24]), 
                          .S3(result_QKT_0[47:36]), 
                          .S4(result_QKT_0[59:48]), 
                          .S5(result_QKT_0[71:60]), 
                          .S6(result_QKT_0[83:72]), 
                          .S7(result_QKT_0[95:84]), 
                          .S8(result_QKT_0[107:96]), 
                          .S9(result_QKT_0[119:108]), 
                          .S10(result_QKT_0[131:120]), 
                          .S11(result_QKT_0[143:132]), 
                          .S12(result_QKT_0[155:144]), 
                          .S13(result_QKT_0[167:156]), 
                          .S14(result_QKT_0[179:168]), 
                          .S15(result_QKT_0[191:180])
                        );

dimc_macro i_dimc_macro_33(.clk(clk_i),
                          .WL(WL_QKT_1), 
                          .wdata(wdata_QKT_1), 
                          .ai(ai_QKT_1), 
                          .RE_(RE_QKT__1), 
                          .PREC(PREC_QKT_1),
                          .PREC_(PREC_QKT__1),
                          .S0(result_QKT_1[11:0]), 
                          .S1(result_QKT_1[23:12]), 
                          .S2(result_QKT_1[35:24]), 
                          .S3(result_QKT_1[47:36]), 
                          .S4(result_QKT_1[59:48]), 
                          .S5(result_QKT_1[71:60]), 
                          .S6(result_QKT_1[83:72]), 
                          .S7(result_QKT_1[95:84]), 
                          .S8(result_QKT_1[107:96]), 
                          .S9(result_QKT_1[119:108]), 
                          .S10(result_QKT_1[131:120]), 
                          .S11(result_QKT_1[143:132]), 
                          .S12(result_QKT_1[155:144]), 
                          .S13(result_QKT_1[167:156]), 
                          .S14(result_QKT_1[179:168]), 
                          .S15(result_QKT_1[191:180])
                        );

dimc_macro i_dimc_macro_34(.clk(clk_i),
                          .WL(WL_QKT_2), 
                          .wdata(wdata_QKT_2), 
                          .ai(ai_QKT_2), 
                          .RE_(RE_QKT__2), 
                          .PREC(PREC_QKT_2),
                          .PREC_(PREC_QKT__2),
                          .S0(result_QKT_2[11:0]), 
                          .S1(result_QKT_2[23:12]), 
                          .S2(result_QKT_2[35:24]), 
                          .S3(result_QKT_2[47:36]), 
                          .S4(result_QKT_2[59:48]), 
                          .S5(result_QKT_2[71:60]), 
                          .S6(result_QKT_2[83:72]), 
                          .S7(result_QKT_2[95:84]), 
                          .S8(result_QKT_2[107:96]), 
                          .S9(result_QKT_2[119:108]), 
                          .S10(result_QKT_2[131:120]), 
                          .S11(result_QKT_2[143:132]), 
                          .S12(result_QKT_2[155:144]), 
                          .S13(result_QKT_2[167:156]), 
                          .S14(result_QKT_2[179:168]), 
                          .S15(result_QKT_2[191:180])
                        );

dimc_macro i_dimc_macro_35(.clk(clk_i),
                          .WL(WL_QKT_3), 
                          .wdata(wdata_QKT_3), 
                          .ai(ai_QKT_3), 
                          .RE_(RE_QKT__3), 
                          .PREC(PREC_QKT_3),
                          .PREC_(PREC_QKT__3),
                          .S0(result_QKT_3[11:0]), 
                          .S1(result_QKT_3[23:12]), 
                          .S2(result_QKT_3[35:24]), 
                          .S3(result_QKT_3[47:36]), 
                          .S4(result_QKT_3[59:48]), 
                          .S5(result_QKT_3[71:60]), 
                          .S6(result_QKT_3[83:72]), 
                          .S7(result_QKT_3[95:84]), 
                          .S8(result_QKT_3[107:96]), 
                          .S9(result_QKT_3[119:108]), 
                          .S10(result_QKT_3[131:120]), 
                          .S11(result_QKT_3[143:132]), 
                          .S12(result_QKT_3[155:144]), 
                          .S13(result_QKT_3[167:156]), 
                          .S14(result_QKT_3[179:168]), 
                          .S15(result_QKT_3[191:180])
                        );

`else
dimc_macro i_dimc_macro_0(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_0), 
                          .wdata(wdata_QKV_0), 
                          .ai(ai_QKV_0), 
                          .RE_(RE_QKV__0), 
                          .PREC(PREC_QKV_0),
                          .PREC_(PREC_QKV__0),
                          .S0(result_QKV_0[11:0]), 
                          .S1(result_QKV_0[23:12]), 
                          .S2(result_QKV_0[35:24]), 
                          .S3(result_QKV_0[47:36]), 
                          .S4(result_QKV_0[59:48]), 
                          .S5(result_QKV_0[71:60]), 
                          .S6(result_QKV_0[83:72]), 
                          .S7(result_QKV_0[95:84]), 
                          .S8(result_QKV_0[107:96]), 
                          .S9(result_QKV_0[119:108]), 
                          .S10(result_QKV_0[131:120]), 
                          .S11(result_QKV_0[143:132]), 
                          .S12(result_QKV_0[155:144]), 
                          .S13(result_QKV_0[167:156]), 
                          .S14(result_QKV_0[179:168]), 
                          .S15(result_QKV_0[191:180])
                        );

dimc_macro i_dimc_macro_1(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_1), 
                          .wdata(wdata_QKV_1), 
                          .ai(ai_QKV_1), 
                          .RE_(RE_QKV__1), 
                          .PREC(PREC_QKV_1),
                          .PREC_(PREC_QKV__1),
                          .S0(result_QKV_1[11:0]), 
                          .S1(result_QKV_1[23:12]), 
                          .S2(result_QKV_1[35:24]), 
                          .S3(result_QKV_1[47:36]), 
                          .S4(result_QKV_1[59:48]), 
                          .S5(result_QKV_1[71:60]), 
                          .S6(result_QKV_1[83:72]), 
                          .S7(result_QKV_1[95:84]), 
                          .S8(result_QKV_1[107:96]), 
                          .S9(result_QKV_1[119:108]), 
                          .S10(result_QKV_1[131:120]), 
                          .S11(result_QKV_1[143:132]), 
                          .S12(result_QKV_1[155:144]), 
                          .S13(result_QKV_1[167:156]), 
                          .S14(result_QKV_1[179:168]), 
                          .S15(result_QKV_1[191:180])
                        );

dimc_macro i_dimc_macro_2(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_2), 
                          .wdata(wdata_QKV_2), 
                          .ai(ai_QKV_2), 
                          .RE_(RE_QKV__2), 
                          .PREC(PREC_QKV_2),
                          .PREC_(PREC_QKV__2),
                          .S0(result_QKV_2[11:0]), 
                          .S1(result_QKV_2[23:12]), 
                          .S2(result_QKV_2[35:24]), 
                          .S3(result_QKV_2[47:36]), 
                          .S4(result_QKV_2[59:48]), 
                          .S5(result_QKV_2[71:60]), 
                          .S6(result_QKV_2[83:72]), 
                          .S7(result_QKV_2[95:84]), 
                          .S8(result_QKV_2[107:96]), 
                          .S9(result_QKV_2[119:108]), 
                          .S10(result_QKV_2[131:120]), 
                          .S11(result_QKV_2[143:132]), 
                          .S12(result_QKV_2[155:144]), 
                          .S13(result_QKV_2[167:156]), 
                          .S14(result_QKV_2[179:168]), 
                          .S15(result_QKV_2[191:180])
                        );

dimc_macro i_dimc_macro_3(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_3), 
                          .wdata(wdata_QKV_3), 
                          .ai(ai_QKV_3), 
                          .RE_(RE_QKV__3), 
                          .PREC(PREC_QKV_3),
                          .PREC_(PREC_QKV__3),
                          .S0(result_QKV_3[11:0]),
                          .S1(result_QKV_3[23:12]),
                          .S2(result_QKV_3[35:24]),
                          .S3(result_QKV_3[47:36]),
                          .S4(result_QKV_3[59:48]),
                          .S5(result_QKV_3[71:60]),
                          .S6(result_QKV_3[83:72]),
                          .S7(result_QKV_3[95:84]),
                          .S8(result_QKV_3[107:96]),
                          .S9(result_QKV_3[119:108]),
                          .S10(result_QKV_3[131:120]),
                          .S11(result_QKV_3[143:132]),
                          .S12(result_QKV_3[155:144]),
                          .S13(result_QKV_3[167:156]),
                          .S14(result_QKV_3[179:168]),
                          .S15(result_QKV_3[191:180])
                        );

dimc_macro i_dimc_macro_4(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_4), 
                          .wdata(wdata_QKV_4), 
                          .ai(ai_QKV_4), 
                          .RE_(RE_QKV__4), 
                          .PREC(PREC_QKV_4),
                          .PREC_(PREC_QKV__4),
                          .S0(result_QKV_4[11:0]), 
                          .S1(result_QKV_4[23:12]), 
                          .S2(result_QKV_4[35:24]), 
                          .S3(result_QKV_4[47:36]), 
                          .S4(result_QKV_4[59:48]), 
                          .S5(result_QKV_4[71:60]), 
                          .S6(result_QKV_4[83:72]), 
                          .S7(result_QKV_4[95:84]), 
                          .S8(result_QKV_4[107:96]), 
                          .S9(result_QKV_4[119:108]), 
                          .S10(result_QKV_4[131:120]), 
                          .S11(result_QKV_4[143:132]), 
                          .S12(result_QKV_4[155:144]), 
                          .S13(result_QKV_4[167:156]), 
                          .S14(result_QKV_4[179:168]), 
                          .S15(result_QKV_4[191:180])
                        );

dimc_macro i_dimc_macro_5(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_5), 
                          .wdata(wdata_QKV_5), 
                          .ai(ai_QKV_5), 
                          .RE_(RE_QKV__5), 
                          .PREC(PREC_QKV_5),
                          .PREC_(PREC_QKV__5),
                          .S0(result_QKV_5[11:0]), 
                          .S1(result_QKV_5[23:12]), 
                          .S2(result_QKV_5[35:24]), 
                          .S3(result_QKV_5[47:36]), 
                          .S4(result_QKV_5[59:48]), 
                          .S5(result_QKV_5[71:60]), 
                          .S6(result_QKV_5[83:72]), 
                          .S7(result_QKV_5[95:84]), 
                          .S8(result_QKV_5[107:96]), 
                          .S9(result_QKV_5[119:108]), 
                          .S10(result_QKV_5[131:120]), 
                          .S11(result_QKV_5[143:132]), 
                          .S12(result_QKV_5[155:144]), 
                          .S13(result_QKV_5[167:156]), 
                          .S14(result_QKV_5[179:168]), 
                          .S15(result_QKV_5[191:180])
                        );

dimc_macro i_dimc_macro_6(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_6), 
                          .wdata(wdata_QKV_6), 
                          .ai(ai_QKV_6), 
                          .RE_(RE_QKV__6), 
                          .PREC(PREC_QKV_6),
                          .PREC_(PREC_QKV__6),
                          .S0(result_QKV_6[11:0]), 
                          .S1(result_QKV_6[23:12]), 
                          .S2(result_QKV_6[35:24]), 
                          .S3(result_QKV_6[47:36]), 
                          .S4(result_QKV_6[59:48]), 
                          .S5(result_QKV_6[71:60]), 
                          .S6(result_QKV_6[83:72]), 
                          .S7(result_QKV_6[95:84]), 
                          .S8(result_QKV_6[107:96]), 
                          .S9(result_QKV_6[119:108]), 
                          .S10(result_QKV_6[131:120]), 
                          .S11(result_QKV_6[143:132]), 
                          .S12(result_QKV_6[155:144]), 
                          .S13(result_QKV_6[167:156]), 
                          .S14(result_QKV_6[179:168]), 
                          .S15(result_QKV_6[191:180])
                        );

dimc_macro i_dimc_macro_7(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_7), 
                          .wdata(wdata_QKV_7), 
                          .ai(ai_QKV_7), 
                          .RE_(RE_QKV__7), 
                          .PREC(PREC_QKV_7),
                          .PREC_(PREC_QKV__7),
                          .S0(result_QKV_7[11:0]), 
                          .S1(result_QKV_7[23:12]), 
                          .S2(result_QKV_7[35:24]), 
                          .S3(result_QKV_7[47:36]), 
                          .S4(result_QKV_7[59:48]), 
                          .S5(result_QKV_7[71:60]), 
                          .S6(result_QKV_7[83:72]), 
                          .S7(result_QKV_7[95:84]), 
                          .S8(result_QKV_7[107:96]), 
                          .S9(result_QKV_7[119:108]), 
                          .S10(result_QKV_7[131:120]), 
                          .S11(result_QKV_7[143:132]), 
                          .S12(result_QKV_7[155:144]), 
                          .S13(result_QKV_7[167:156]), 
                          .S14(result_QKV_7[179:168]), 
                          .S15(result_QKV_7[191:180])
                        );

dimc_macro i_dimc_macro_8(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_8), 
                          .wdata(wdata_QKV_8), 
                          .ai(ai_QKV_8), 
                          .RE_(RE_QKV__8), 
                          .PREC(PREC_QKV_8),
                          .PREC_(PREC_QKV__8),
                          .S0(result_QKV_8[11:0]), 
                          .S1(result_QKV_8[23:12]), 
                          .S2(result_QKV_8[35:24]), 
                          .S3(result_QKV_8[47:36]), 
                          .S4(result_QKV_8[59:48]), 
                          .S5(result_QKV_8[71:60]), 
                          .S6(result_QKV_8[83:72]), 
                          .S7(result_QKV_8[95:84]), 
                          .S8(result_QKV_8[107:96]), 
                          .S9(result_QKV_8[119:108]), 
                          .S10(result_QKV_8[131:120]), 
                          .S11(result_QKV_8[143:132]), 
                          .S12(result_QKV_8[155:144]), 
                          .S13(result_QKV_8[167:156]), 
                          .S14(result_QKV_8[179:168]), 
                          .S15(result_QKV_8[191:180])
                        );

dimc_macro i_dimc_macro_9(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_9), 
                          .wdata(wdata_QKV_9), 
                          .ai(ai_QKV_9), 
                          .RE_(RE_QKV__9), 
                          .PREC(PREC_QKV_9),
                          .PREC_(PREC_QKV__9),
                          .S0(result_QKV_9[11:0]), 
                          .S1(result_QKV_9[23:12]), 
                          .S2(result_QKV_9[35:24]), 
                          .S3(result_QKV_9[47:36]), 
                          .S4(result_QKV_9[59:48]), 
                          .S5(result_QKV_9[71:60]), 
                          .S6(result_QKV_9[83:72]), 
                          .S7(result_QKV_9[95:84]), 
                          .S8(result_QKV_9[107:96]), 
                          .S9(result_QKV_9[119:108]), 
                          .S10(result_QKV_9[131:120]), 
                          .S11(result_QKV_9[143:132]), 
                          .S12(result_QKV_9[155:144]), 
                          .S13(result_QKV_9[167:156]), 
                          .S14(result_QKV_9[179:168]), 
                          .S15(result_QKV_9[191:180])
                        );

dimc_macro i_dimc_macro_10(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_10), 
                          .wdata(wdata_QKV_10), 
                          .ai(ai_QKV_10), 
                          .RE_(RE_QKV__10), 
                          .PREC(PREC_QKV_10),
                          .PREC_(PREC_QKV__10),
                          .S0(result_QKV_10[11:0]), 
                          .S1(result_QKV_10[23:12]), 
                          .S2(result_QKV_10[35:24]), 
                          .S3(result_QKV_10[47:36]), 
                          .S4(result_QKV_10[59:48]), 
                          .S5(result_QKV_10[71:60]), 
                          .S6(result_QKV_10[83:72]), 
                          .S7(result_QKV_10[95:84]), 
                          .S8(result_QKV_10[107:96]), 
                          .S9(result_QKV_10[119:108]), 
                          .S10(result_QKV_10[131:120]), 
                          .S11(result_QKV_10[143:132]), 
                          .S12(result_QKV_10[155:144]), 
                          .S13(result_QKV_10[167:156]), 
                          .S14(result_QKV_10[179:168]), 
                          .S15(result_QKV_10[191:180])
                        );

dimc_macro i_dimc_macro_11(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_11), 
                          .wdata(wdata_QKV_11), 
                          .ai(ai_QKV_11), 
                          .RE_(RE_QKV__11), 
                          .PREC(PREC_QKV_11),
                          .PREC_(PREC_QKV__11),
                          .S0(result_QKV_11[11:0]), 
                          .S1(result_QKV_11[23:12]), 
                          .S2(result_QKV_11[35:24]), 
                          .S3(result_QKV_11[47:36]), 
                          .S4(result_QKV_11[59:48]), 
                          .S5(result_QKV_11[71:60]), 
                          .S6(result_QKV_11[83:72]), 
                          .S7(result_QKV_11[95:84]), 
                          .S8(result_QKV_11[107:96]), 
                          .S9(result_QKV_11[119:108]), 
                          .S10(result_QKV_11[131:120]), 
                          .S11(result_QKV_11[143:132]), 
                          .S12(result_QKV_11[155:144]), 
                          .S13(result_QKV_11[167:156]), 
                          .S14(result_QKV_11[179:168]), 
                          .S15(result_QKV_11[191:180])
                        );

dimc_macro i_dimc_macro_12(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_12), 
                          .wdata(wdata_QKV_12), 
                          .ai(ai_QKV_12), 
                          .RE_(RE_QKV__12), 
                          .PREC(PREC_QKV_12),
                          .PREC_(PREC_QKV__12),
                          .S0(result_QKV_12[11:0]), 
                          .S1(result_QKV_12[23:12]), 
                          .S2(result_QKV_12[35:24]), 
                          .S3(result_QKV_12[47:36]), 
                          .S4(result_QKV_12[59:48]), 
                          .S5(result_QKV_12[71:60]), 
                          .S6(result_QKV_12[83:72]), 
                          .S7(result_QKV_12[95:84]), 
                          .S8(result_QKV_12[107:96]), 
                          .S9(result_QKV_12[119:108]), 
                          .S10(result_QKV_12[131:120]), 
                          .S11(result_QKV_12[143:132]), 
                          .S12(result_QKV_12[155:144]), 
                          .S13(result_QKV_12[167:156]), 
                          .S14(result_QKV_12[179:168]), 
                          .S15(result_QKV_12[191:180])
                        );

dimc_macro i_dimc_macro_13(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_13), 
                          .wdata(wdata_QKV_13), 
                          .ai(ai_QKV_13), 
                          .RE_(RE_QKV__13), 
                          .PREC(PREC_QKV_13),
                          .PREC_(PREC_QKV__13),
                          .S0(result_QKV_13[11:0]), 
                          .S1(result_QKV_13[23:12]), 
                          .S2(result_QKV_13[35:24]), 
                          .S3(result_QKV_13[47:36]), 
                          .S4(result_QKV_13[59:48]), 
                          .S5(result_QKV_13[71:60]), 
                          .S6(result_QKV_13[83:72]), 
                          .S7(result_QKV_13[95:84]), 
                          .S8(result_QKV_13[107:96]), 
                          .S9(result_QKV_13[119:108]), 
                          .S10(result_QKV_13[131:120]), 
                          .S11(result_QKV_13[143:132]), 
                          .S12(result_QKV_13[155:144]), 
                          .S13(result_QKV_13[167:156]), 
                          .S14(result_QKV_13[179:168]), 
                          .S15(result_QKV_13[191:180])
                        );

dimc_macro i_dimc_macro_14(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_14), 
                          .wdata(wdata_QKV_14), 
                          .ai(ai_QKV_14), 
                          .RE_(RE_QKV__14), 
                          .PREC(PREC_QKV_14),
                          .PREC_(PREC_QKV__14),
                          .S0(result_QKV_14[11:0]), 
                          .S1(result_QKV_14[23:12]), 
                          .S2(result_QKV_14[35:24]), 
                          .S3(result_QKV_14[47:36]), 
                          .S4(result_QKV_14[59:48]), 
                          .S5(result_QKV_14[71:60]), 
                          .S6(result_QKV_14[83:72]), 
                          .S7(result_QKV_14[95:84]), 
                          .S8(result_QKV_14[107:96]), 
                          .S9(result_QKV_14[119:108]), 
                          .S10(result_QKV_14[131:120]), 
                          .S11(result_QKV_14[143:132]), 
                          .S12(result_QKV_14[155:144]), 
                          .S13(result_QKV_14[167:156]), 
                          .S14(result_QKV_14[179:168]), 
                          .S15(result_QKV_14[191:180])
                        );

dimc_macro i_dimc_macro_15(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_15), 
                          .wdata(wdata_QKV_15), 
                          .ai(ai_QKV_15), 
                          .RE_(RE_QKV__15), 
                          .PREC(PREC_QKV_15),
                          .PREC_(PREC_QKV__15),
                          .S0(result_QKV_15[11:0]), 
                          .S1(result_QKV_15[23:12]), 
                          .S2(result_QKV_15[35:24]), 
                          .S3(result_QKV_15[47:36]), 
                          .S4(result_QKV_15[59:48]), 
                          .S5(result_QKV_15[71:60]), 
                          .S6(result_QKV_15[83:72]), 
                          .S7(result_QKV_15[95:84]), 
                          .S8(result_QKV_15[107:96]), 
                          .S9(result_QKV_15[119:108]), 
                          .S10(result_QKV_15[131:120]), 
                          .S11(result_QKV_15[143:132]), 
                          .S12(result_QKV_15[155:144]), 
                          .S13(result_QKV_15[167:156]), 
                          .S14(result_QKV_15[179:168]), 
                          .S15(result_QKV_15[191:180])
                        );

dimc_macro i_dimc_macro_16(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_16), 
                          .wdata(wdata_QKV_16), 
                          .ai(ai_QKV_16), 
                          .RE_(RE_QKV__16), 
                          .PREC(PREC_QKV_16),
                          .PREC_(PREC_QKV__16),
                          .S0(result_QKV_16[11:0]), 
                          .S1(result_QKV_16[23:12]), 
                          .S2(result_QKV_16[35:24]), 
                          .S3(result_QKV_16[47:36]), 
                          .S4(result_QKV_16[59:48]), 
                          .S5(result_QKV_16[71:60]), 
                          .S6(result_QKV_16[83:72]), 
                          .S7(result_QKV_16[95:84]), 
                          .S8(result_QKV_16[107:96]), 
                          .S9(result_QKV_16[119:108]), 
                          .S10(result_QKV_16[131:120]), 
                          .S11(result_QKV_16[143:132]), 
                          .S12(result_QKV_16[155:144]), 
                          .S13(result_QKV_16[167:156]), 
                          .S14(result_QKV_16[179:168]), 
                          .S15(result_QKV_16[191:180])
                        );

dimc_macro i_dimc_macro_17(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_17), 
                          .wdata(wdata_QKV_17), 
                          .ai(ai_QKV_17), 
                          .RE_(RE_QKV__17), 
                          .PREC(PREC_QKV_17),
                          .PREC_(PREC_QKV__17),
                          .S0(result_QKV_17[11:0]), 
                          .S1(result_QKV_17[23:12]), 
                          .S2(result_QKV_17[35:24]), 
                          .S3(result_QKV_17[47:36]), 
                          .S4(result_QKV_17[59:48]), 
                          .S5(result_QKV_17[71:60]), 
                          .S6(result_QKV_17[83:72]), 
                          .S7(result_QKV_17[95:84]), 
                          .S8(result_QKV_17[107:96]), 
                          .S9(result_QKV_17[119:108]), 
                          .S10(result_QKV_17[131:120]), 
                          .S11(result_QKV_17[143:132]), 
                          .S12(result_QKV_17[155:144]), 
                          .S13(result_QKV_17[167:156]), 
                          .S14(result_QKV_17[179:168]), 
                          .S15(result_QKV_17[191:180])
                        );

dimc_macro i_dimc_macro_18(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_18), 
                          .wdata(wdata_QKV_18), 
                          .ai(ai_QKV_18), 
                          .RE_(RE_QKV__18), 
                          .PREC(PREC_QKV_18),
                          .PREC_(PREC_QKV__18),
                          .S0(result_QKV_18[11:0]), 
                          .S1(result_QKV_18[23:12]), 
                          .S2(result_QKV_18[35:24]), 
                          .S3(result_QKV_18[47:36]), 
                          .S4(result_QKV_18[59:48]), 
                          .S5(result_QKV_18[71:60]), 
                          .S6(result_QKV_18[83:72]), 
                          .S7(result_QKV_18[95:84]), 
                          .S8(result_QKV_18[107:96]), 
                          .S9(result_QKV_18[119:108]), 
                          .S10(result_QKV_18[131:120]), 
                          .S11(result_QKV_18[143:132]), 
                          .S12(result_QKV_18[155:144]), 
                          .S13(result_QKV_18[167:156]), 
                          .S14(result_QKV_18[179:168]), 
                          .S15(result_QKV_18[191:180])
                        );

dimc_macro i_dimc_macro_19(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_19), 
                          .wdata(wdata_QKV_19), 
                          .ai(ai_QKV_19), 
                          .RE_(RE_QKV__19), 
                          .PREC(PREC_QKV_19),
                          .PREC_(PREC_QKV__19),
                          .S0(result_QKV_19[11:0]), 
                          .S1(result_QKV_19[23:12]), 
                          .S2(result_QKV_19[35:24]), 
                          .S3(result_QKV_19[47:36]), 
                          .S4(result_QKV_19[59:48]), 
                          .S5(result_QKV_19[71:60]), 
                          .S6(result_QKV_19[83:72]), 
                          .S7(result_QKV_19[95:84]), 
                          .S8(result_QKV_19[107:96]), 
                          .S9(result_QKV_19[119:108]), 
                          .S10(result_QKV_19[131:120]), 
                          .S11(result_QKV_19[143:132]), 
                          .S12(result_QKV_19[155:144]), 
                          .S13(result_QKV_19[167:156]), 
                          .S14(result_QKV_19[179:168]), 
                          .S15(result_QKV_19[191:180])
                        );

dimc_macro i_dimc_macro_20(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_20), 
                          .wdata(wdata_QKV_20), 
                          .ai(ai_QKV_20), 
                          .RE_(RE_QKV__20), 
                          .PREC(PREC_QKV_20),
                          .PREC_(PREC_QKV__20),
                          .S0(result_QKV_20[11:0]), 
                          .S1(result_QKV_20[23:12]), 
                          .S2(result_QKV_20[35:24]), 
                          .S3(result_QKV_20[47:36]), 
                          .S4(result_QKV_20[59:48]), 
                          .S5(result_QKV_20[71:60]), 
                          .S6(result_QKV_20[83:72]), 
                          .S7(result_QKV_20[95:84]), 
                          .S8(result_QKV_20[107:96]), 
                          .S9(result_QKV_20[119:108]), 
                          .S10(result_QKV_20[131:120]), 
                          .S11(result_QKV_20[143:132]), 
                          .S12(result_QKV_20[155:144]), 
                          .S13(result_QKV_20[167:156]), 
                          .S14(result_QKV_20[179:168]), 
                          .S15(result_QKV_20[191:180])
                        );

dimc_macro i_dimc_macro_21(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_21), 
                          .wdata(wdata_QKV_21), 
                          .ai(ai_QKV_21), 
                          .RE_(RE_QKV__21), 
                          .PREC(PREC_QKV_21),
                          .PREC_(PREC_QKV__21),
                          .S0(result_QKV_21[11:0]), 
                          .S1(result_QKV_21[23:12]), 
                          .S2(result_QKV_21[35:24]), 
                          .S3(result_QKV_21[47:36]), 
                          .S4(result_QKV_21[59:48]), 
                          .S5(result_QKV_21[71:60]), 
                          .S6(result_QKV_21[83:72]), 
                          .S7(result_QKV_21[95:84]), 
                          .S8(result_QKV_21[107:96]), 
                          .S9(result_QKV_21[119:108]), 
                          .S10(result_QKV_21[131:120]), 
                          .S11(result_QKV_21[143:132]), 
                          .S12(result_QKV_21[155:144]), 
                          .S13(result_QKV_21[167:156]), 
                          .S14(result_QKV_21[179:168]), 
                          .S15(result_QKV_21[191:180])
                        );

dimc_macro i_dimc_macro_22(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_22), 
                          .wdata(wdata_QKV_22), 
                          .ai(ai_QKV_22), 
                          .RE_(RE_QKV__22), 
                          .PREC(PREC_QKV_22),
                          .PREC_(PREC_QKV__22),
                          .S0(result_QKV_22[11:0]), 
                          .S1(result_QKV_22[23:12]), 
                          .S2(result_QKV_22[35:24]), 
                          .S3(result_QKV_22[47:36]), 
                          .S4(result_QKV_22[59:48]), 
                          .S5(result_QKV_22[71:60]), 
                          .S6(result_QKV_22[83:72]), 
                          .S7(result_QKV_22[95:84]), 
                          .S8(result_QKV_22[107:96]), 
                          .S9(result_QKV_22[119:108]), 
                          .S10(result_QKV_22[131:120]), 
                          .S11(result_QKV_22[143:132]), 
                          .S12(result_QKV_22[155:144]), 
                          .S13(result_QKV_22[167:156]), 
                          .S14(result_QKV_22[179:168]), 
                          .S15(result_QKV_22[191:180])
                        );

dimc_macro i_dimc_macro_23(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_23), 
                          .wdata(wdata_QKV_23), 
                          .ai(ai_QKV_23), 
                          .RE_(RE_QKV__23), 
                          .PREC(PREC_QKV_23),
                          .PREC_(PREC_QKV__23),
                          .S0(result_QKV_23[11:0]), 
                          .S1(result_QKV_23[23:12]), 
                          .S2(result_QKV_23[35:24]), 
                          .S3(result_QKV_23[47:36]), 
                          .S4(result_QKV_23[59:48]), 
                          .S5(result_QKV_23[71:60]), 
                          .S6(result_QKV_23[83:72]), 
                          .S7(result_QKV_23[95:84]), 
                          .S8(result_QKV_23[107:96]), 
                          .S9(result_QKV_23[119:108]), 
                          .S10(result_QKV_23[131:120]), 
                          .S11(result_QKV_23[143:132]), 
                          .S12(result_QKV_23[155:144]), 
                          .S13(result_QKV_23[167:156]), 
                          .S14(result_QKV_23[179:168]), 
                          .S15(result_QKV_23[191:180])
                        );

dimc_macro i_dimc_macro_24(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_24), 
                          .wdata(wdata_QKV_24), 
                          .ai(ai_QKV_24), 
                          .RE_(RE_QKV__24), 
                          .PREC(PREC_QKV_24),
                          .PREC_(PREC_QKV__24),
                          .S0(result_QKV_24[11:0]), 
                          .S1(result_QKV_24[23:12]), 
                          .S2(result_QKV_24[35:24]), 
                          .S3(result_QKV_24[47:36]), 
                          .S4(result_QKV_24[59:48]), 
                          .S5(result_QKV_24[71:60]), 
                          .S6(result_QKV_24[83:72]), 
                          .S7(result_QKV_24[95:84]), 
                          .S8(result_QKV_24[107:96]), 
                          .S9(result_QKV_24[119:108]), 
                          .S10(result_QKV_24[131:120]), 
                          .S11(result_QKV_24[143:132]), 
                          .S12(result_QKV_24[155:144]), 
                          .S13(result_QKV_24[167:156]), 
                          .S14(result_QKV_24[179:168]), 
                          .S15(result_QKV_24[191:180])
                        );

dimc_macro i_dimc_macro_25(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_25), 
                          .wdata(wdata_QKV_25), 
                          .ai(ai_QKV_25), 
                          .RE_(RE_QKV__25), 
                          .PREC(PREC_QKV_25),
                          .PREC_(PREC_QKV__25),
                          .S0(result_QKV_25[11:0]), 
                          .S1(result_QKV_25[23:12]), 
                          .S2(result_QKV_25[35:24]), 
                          .S3(result_QKV_25[47:36]), 
                          .S4(result_QKV_25[59:48]), 
                          .S5(result_QKV_25[71:60]), 
                          .S6(result_QKV_25[83:72]), 
                          .S7(result_QKV_25[95:84]), 
                          .S8(result_QKV_25[107:96]), 
                          .S9(result_QKV_25[119:108]), 
                          .S10(result_QKV_25[131:120]), 
                          .S11(result_QKV_25[143:132]), 
                          .S12(result_QKV_25[155:144]), 
                          .S13(result_QKV_25[167:156]), 
                          .S14(result_QKV_25[179:168]), 
                          .S15(result_QKV_25[191:180])
                        );

dimc_macro i_dimc_macro_26(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_26), 
                          .wdata(wdata_QKV_26), 
                          .ai(ai_QKV_26), 
                          .RE_(RE_QKV__26), 
                          .PREC(PREC_QKV_26),
                          .PREC_(PREC_QKV__26),
                          .S0(result_QKV_26[11:0]), 
                          .S1(result_QKV_26[23:12]), 
                          .S2(result_QKV_26[35:24]), 
                          .S3(result_QKV_26[47:36]), 
                          .S4(result_QKV_26[59:48]), 
                          .S5(result_QKV_26[71:60]), 
                          .S6(result_QKV_26[83:72]), 
                          .S7(result_QKV_26[95:84]), 
                          .S8(result_QKV_26[107:96]), 
                          .S9(result_QKV_26[119:108]), 
                          .S10(result_QKV_26[131:120]), 
                          .S11(result_QKV_26[143:132]), 
                          .S12(result_QKV_26[155:144]), 
                          .S13(result_QKV_26[167:156]), 
                          .S14(result_QKV_26[179:168]), 
                          .S15(result_QKV_26[191:180])
                        );

dimc_macro i_dimc_macro_27(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_27), 
                          .wdata(wdata_QKV_27), 
                          .ai(ai_QKV_27), 
                          .RE_(RE_QKV__27), 
                          .PREC(PREC_QKV_27),
                          .PREC_(PREC_QKV__27),
                          .S0(result_QKV_27[11:0]), 
                          .S1(result_QKV_27[23:12]), 
                          .S2(result_QKV_27[35:24]), 
                          .S3(result_QKV_27[47:36]), 
                          .S4(result_QKV_27[59:48]), 
                          .S5(result_QKV_27[71:60]), 
                          .S6(result_QKV_27[83:72]), 
                          .S7(result_QKV_27[95:84]), 
                          .S8(result_QKV_27[107:96]), 
                          .S9(result_QKV_27[119:108]), 
                          .S10(result_QKV_27[131:120]), 
                          .S11(result_QKV_27[143:132]), 
                          .S12(result_QKV_27[155:144]), 
                          .S13(result_QKV_27[167:156]), 
                          .S14(result_QKV_27[179:168]), 
                          .S15(result_QKV_27[191:180])
                        );

dimc_macro i_dimc_macro_28(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_28), 
                          .wdata(wdata_QKV_28), 
                          .ai(ai_QKV_28), 
                          .RE_(RE_QKV__28), 
                          .PREC(PREC_QKV_28),
                          .PREC_(PREC_QKV__28),
                          .S0(result_QKV_28[11:0]), 
                          .S1(result_QKV_28[23:12]), 
                          .S2(result_QKV_28[35:24]), 
                          .S3(result_QKV_28[47:36]), 
                          .S4(result_QKV_28[59:48]), 
                          .S5(result_QKV_28[71:60]), 
                          .S6(result_QKV_28[83:72]), 
                          .S7(result_QKV_28[95:84]), 
                          .S8(result_QKV_28[107:96]), 
                          .S9(result_QKV_28[119:108]), 
                          .S10(result_QKV_28[131:120]), 
                          .S11(result_QKV_28[143:132]), 
                          .S12(result_QKV_28[155:144]), 
                          .S13(result_QKV_28[167:156]), 
                          .S14(result_QKV_28[179:168]), 
                          .S15(result_QKV_28[191:180])
                        );

dimc_macro i_dimc_macro_29(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_29), 
                          .wdata(wdata_QKV_29), 
                          .ai(ai_QKV_29), 
                          .RE_(RE_QKV__29), 
                          .PREC(PREC_QKV_29),
                          .PREC_(PREC_QKV__29),
                          .S0(result_QKV_29[11:0]), 
                          .S1(result_QKV_29[23:12]), 
                          .S2(result_QKV_29[35:24]), 
                          .S3(result_QKV_29[47:36]), 
                          .S4(result_QKV_29[59:48]), 
                          .S5(result_QKV_29[71:60]), 
                          .S6(result_QKV_29[83:72]), 
                          .S7(result_QKV_29[95:84]), 
                          .S8(result_QKV_29[107:96]), 
                          .S9(result_QKV_29[119:108]), 
                          .S10(result_QKV_29[131:120]), 
                          .S11(result_QKV_29[143:132]), 
                          .S12(result_QKV_29[155:144]), 
                          .S13(result_QKV_29[167:156]), 
                          .S14(result_QKV_29[179:168]), 
                          .S15(result_QKV_29[191:180])
                        );

dimc_macro i_dimc_macro_30(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_30), 
                          .wdata(wdata_QKV_30), 
                          .ai(ai_QKV_30), 
                          .RE_(RE_QKV__30), 
                          .PREC(PREC_QKV_30),
                          .PREC_(PREC_QKV__30),
                          .S0(result_QKV_30[11:0]), 
                          .S1(result_QKV_30[23:12]), 
                          .S2(result_QKV_30[35:24]), 
                          .S3(result_QKV_30[47:36]), 
                          .S4(result_QKV_30[59:48]), 
                          .S5(result_QKV_30[71:60]), 
                          .S6(result_QKV_30[83:72]), 
                          .S7(result_QKV_30[95:84]), 
                          .S8(result_QKV_30[107:96]), 
                          .S9(result_QKV_30[119:108]), 
                          .S10(result_QKV_30[131:120]), 
                          .S11(result_QKV_30[143:132]), 
                          .S12(result_QKV_30[155:144]), 
                          .S13(result_QKV_30[167:156]), 
                          .S14(result_QKV_30[179:168]), 
                          .S15(result_QKV_30[191:180])
                        );

dimc_macro i_dimc_macro_31(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKV_31), 
                          .wdata(wdata_QKV_31), 
                          .ai(ai_QKV_31), 
                          .RE_(RE_QKV__31), 
                          .PREC(PREC_QKV_31),
                          .PREC_(PREC_QKV__31),
                          .S0(result_QKV_31[11:0]), 
                          .S1(result_QKV_31[23:12]), 
                          .S2(result_QKV_31[35:24]), 
                          .S3(result_QKV_31[47:36]), 
                          .S4(result_QKV_31[59:48]), 
                          .S5(result_QKV_31[71:60]), 
                          .S6(result_QKV_31[83:72]), 
                          .S7(result_QKV_31[95:84]), 
                          .S8(result_QKV_31[107:96]), 
                          .S9(result_QKV_31[119:108]), 
                          .S10(result_QKV_31[131:120]), 
                          .S11(result_QKV_31[143:132]), 
                          .S12(result_QKV_31[155:144]), 
                          .S13(result_QKV_31[167:156]), 
                          .S14(result_QKV_31[179:168]), 
                          .S15(result_QKV_31[191:180])
                        );

dimc_macro i_dimc_macro_32(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKT_0), 
                          .wdata(wdata_QKT_0), 
                          .ai(ai_QKT_0), 
                          .RE_(RE_QKT__0), 
                          .PREC(PREC_QKT_0),
                          .PREC_(PREC_QKT__0),
                          .S0(result_QKT_0[11:0]), 
                          .S1(result_QKT_0[23:12]), 
                          .S2(result_QKT_0[35:24]), 
                          .S3(result_QKT_0[47:36]), 
                          .S4(result_QKT_0[59:48]), 
                          .S5(result_QKT_0[71:60]), 
                          .S6(result_QKT_0[83:72]), 
                          .S7(result_QKT_0[95:84]), 
                          .S8(result_QKT_0[107:96]), 
                          .S9(result_QKT_0[119:108]), 
                          .S10(result_QKT_0[131:120]), 
                          .S11(result_QKT_0[143:132]), 
                          .S12(result_QKT_0[155:144]), 
                          .S13(result_QKT_0[167:156]), 
                          .S14(result_QKT_0[179:168]), 
                          .S15(result_QKT_0[191:180])
                        );

dimc_macro i_dimc_macro_33(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKT_1), 
                          .wdata(wdata_QKT_1), 
                          .ai(ai_QKT_1), 
                          .RE_(RE_QKT__1), 
                          .PREC(PREC_QKT_1),
                          .PREC_(PREC_QKT__1),
                          .S0(result_QKT_1[11:0]), 
                          .S1(result_QKT_1[23:12]), 
                          .S2(result_QKT_1[35:24]), 
                          .S3(result_QKT_1[47:36]), 
                          .S4(result_QKT_1[59:48]), 
                          .S5(result_QKT_1[71:60]), 
                          .S6(result_QKT_1[83:72]), 
                          .S7(result_QKT_1[95:84]), 
                          .S8(result_QKT_1[107:96]), 
                          .S9(result_QKT_1[119:108]), 
                          .S10(result_QKT_1[131:120]), 
                          .S11(result_QKT_1[143:132]), 
                          .S12(result_QKT_1[155:144]), 
                          .S13(result_QKT_1[167:156]), 
                          .S14(result_QKT_1[179:168]), 
                          .S15(result_QKT_1[191:180])
                        );

dimc_macro i_dimc_macro_34(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKT_2), 
                          .wdata(wdata_QKT_2), 
                          .ai(ai_QKT_2), 
                          .RE_(RE_QKT__2), 
                          .PREC(PREC_QKT_2),
                          .PREC_(PREC_QKT__2),
                          .S0(result_QKT_2[11:0]), 
                          .S1(result_QKT_2[23:12]), 
                          .S2(result_QKT_2[35:24]), 
                          .S3(result_QKT_2[47:36]), 
                          .S4(result_QKT_2[59:48]), 
                          .S5(result_QKT_2[71:60]), 
                          .S6(result_QKT_2[83:72]), 
                          .S7(result_QKT_2[95:84]), 
                          .S8(result_QKT_2[107:96]), 
                          .S9(result_QKT_2[119:108]), 
                          .S10(result_QKT_2[131:120]), 
                          .S11(result_QKT_2[143:132]), 
                          .S12(result_QKT_2[155:144]), 
                          .S13(result_QKT_2[167:156]), 
                          .S14(result_QKT_2[179:168]), 
                          .S15(result_QKT_2[191:180])
                        );

dimc_macro i_dimc_macro_35(.clk(clk_i),
                          .rst(rst),
                          .WL(WL_QKT_3), 
                          .wdata(wdata_QKT_3), 
                          .ai(ai_QKT_3), 
                          .RE_(RE_QKT__3), 
                          .PREC(PREC_QKT_3),
                          .PREC_(PREC_QKT__3),
                          .S0(result_QKT_3[11:0]), 
                          .S1(result_QKT_3[23:12]), 
                          .S2(result_QKT_3[35:24]), 
                          .S3(result_QKT_3[47:36]), 
                          .S4(result_QKT_3[59:48]), 
                          .S5(result_QKT_3[71:60]), 
                          .S6(result_QKT_3[83:72]), 
                          .S7(result_QKT_3[95:84]), 
                          .S8(result_QKT_3[107:96]), 
                          .S9(result_QKT_3[119:108]), 
                          .S10(result_QKT_3[131:120]), 
                          .S11(result_QKT_3[143:132]), 
                          .S12(result_QKT_3[155:144]), 
                          .S13(result_QKT_3[167:156]), 
                          .S14(result_QKT_3[179:168]), 
                          .S15(result_QKT_3[191:180])
                        );

`endif

endmodule
