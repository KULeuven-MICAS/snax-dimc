`timescale 1ps / 1ps
module qkt_macro_handler_hub_Div_32Ux32U_8U_4(
          in2,
          in1,
          out1,
          clk,
          stall,
          clr
);
   input [31:0] in2;
   input [31:0] in1;
   output [7:0] out1;
   input clk;
   input stall;
   input clr;
wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13,
     n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25,
     n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37,
     n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49,
     n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61,
     n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73,
     n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85,
     n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97,
     n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108,
     n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119,
     n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130,
     n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141,
     n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152,
     n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163,
     n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174,
     n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185,
     n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196,
     n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207,
     n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218,
     n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229,
     n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240,
     n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251,
     n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262,
     n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273,
     n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284,
     n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295,
     n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306,
     n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317,
     n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328,
     n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339,
     n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350,
     n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361,
     n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372,
     n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383,
     n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394,
     n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405,
     n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416,
     n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427,
     n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438,
     n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449,
     n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460,
     n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471,
     n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482,
     n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493,
     n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504,
     n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515,
     n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526,
     n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537,
     n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548,
     n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559,
     n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570,
     n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581,
     n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592,
     n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603,
     n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614,
     n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625,
     n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636,
     n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646, n_647,
     n_648, n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658,
     n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669,
     n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680,
     n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691,
     n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702,
     n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713,
     n_714, n_715, n_716, n_717, n_718, n_719, n_720, sub_230_64_n_0,
     sub_230_64_n_2, sub_230_64_n_3, sub_230_64_n_4, sub_230_64_n_5,
     sub_230_64_n_6, sub_230_64_n_7, sub_230_64_n_8, sub_230_64_n_9,
     sub_230_64_n_10, sub_230_64_n_11, sub_230_64_n_12, sub_230_64_n_13,
     sub_230_64_n_14, sub_230_64_n_15, sub_230_64_n_16, sub_230_64_n_17,
     sub_230_64_n_18, sub_230_64_n_19, sub_230_64_n_20, sub_230_64_n_22,
     sub_230_64_n_23, sub_230_64_n_24, sub_230_64_n_25, sub_230_64_n_26,
     sub_230_64_n_27, sub_260_63_n_0, sub_260_63_n_1, sub_260_63_n_4,
     sub_260_63_n_5, sub_260_63_n_6, sub_260_63_n_7, sub_260_63_n_8,
     sub_260_63_n_9, sub_260_63_n_10, sub_260_63_n_11, sub_260_63_n_12,
     sub_260_63_n_13, sub_260_63_n_14, sub_260_63_n_15, sub_260_63_n_16,
     sub_260_63_n_17, sub_260_63_n_18, sub_260_63_n_19, sub_260_63_n_20,
     sub_260_63_n_21, sub_260_63_n_22, sub_260_63_n_23, sub_260_63_n_24,
     sub_260_63_n_25, sub_260_63_n_26, sub_260_63_n_28, sub_260_63_n_29,
     sub_260_63_n_30, sub_260_63_n_31, sub_260_63_n_32, sub_260_63_n_33,
     sub_260_63_n_34, sub_260_63_n_35, sub_260_63_n_36, sub_260_63_n_37,
     sub_290_62_n_1, sub_290_62_n_2, sub_290_62_n_3, sub_290_62_n_4,
     sub_290_62_n_5, sub_290_62_n_6, sub_290_62_n_8, sub_290_62_n_9,
     sub_290_62_n_10, sub_290_62_n_11, sub_290_62_n_12, sub_290_62_n_13,
     sub_290_62_n_14, sub_290_62_n_15, sub_290_62_n_16, sub_290_62_n_17,
     sub_290_62_n_18, sub_290_62_n_19, sub_290_62_n_20, sub_290_62_n_21,
     sub_290_62_n_22, sub_290_62_n_23, sub_290_62_n_24, sub_290_62_n_25,
     sub_290_62_n_26, sub_290_62_n_27, sub_290_62_n_28, sub_290_62_n_29,
     sub_290_62_n_30, sub_290_62_n_31, sub_290_62_n_33, sub_290_62_n_34,
     sub_290_62_n_35, sub_290_62_n_36, sub_290_62_n_37, sub_290_62_n_38,
     sub_290_62_n_39, sub_290_62_n_40, sub_320_61_n_0, sub_320_61_n_1,
     sub_320_61_n_2, sub_320_61_n_3, sub_320_61_n_4, sub_320_61_n_6,
     sub_320_61_n_7, sub_320_61_n_8, sub_320_61_n_9, sub_320_61_n_10,
     sub_320_61_n_11, sub_320_61_n_12, sub_320_61_n_13, sub_320_61_n_14,
     sub_320_61_n_15, sub_320_61_n_16, sub_320_61_n_17, sub_320_61_n_18,
     sub_320_61_n_19, sub_320_61_n_20, sub_320_61_n_21, sub_320_61_n_22,
     sub_320_61_n_23, sub_320_61_n_24, sub_320_61_n_25, sub_320_61_n_26,
     sub_320_61_n_27, sub_320_61_n_28, sub_320_61_n_30, sub_320_61_n_31,
     sub_320_61_n_32, sub_320_61_n_33, sub_320_61_n_34, sub_320_61_n_35,
     sub_320_61_n_36, sub_320_61_n_38, sub_320_61_n_39, sub_320_61_n_40,
     sub_320_61_n_41, sub_320_61_n_43, sub_320_61_n_44, sub_320_61_n_45,
     sub_350_60_n_0, sub_350_60_n_1, sub_350_60_n_2, sub_350_60_n_3,
     sub_350_60_n_4, sub_350_60_n_5, sub_350_60_n_7, sub_350_60_n_8,
     sub_350_60_n_9, sub_350_60_n_10, sub_350_60_n_11, sub_350_60_n_12,
     sub_350_60_n_13, sub_350_60_n_14, sub_350_60_n_15, sub_350_60_n_16,
     sub_350_60_n_17, sub_350_60_n_18, sub_350_60_n_19, sub_350_60_n_20,
     sub_350_60_n_21, sub_350_60_n_22, sub_350_60_n_23, sub_350_60_n_24,
     sub_350_60_n_25, sub_350_60_n_26, sub_350_60_n_27, sub_350_60_n_28,
     sub_350_60_n_29, sub_350_60_n_30, sub_350_60_n_31, sub_350_60_n_32,
     sub_350_60_n_33, sub_350_60_n_34, sub_350_60_n_36, sub_350_60_n_37,
     sub_350_60_n_38, sub_350_60_n_39, sub_350_60_n_40, sub_350_60_n_41,
     sub_350_60_n_42, sub_350_60_n_43, sub_350_60_n_44, sub_350_60_n_45,
     sub_350_60_n_46, sub_350_60_n_47, sub_350_60_n_49, sub_350_60_n_50,
     sub_350_60_n_51, sub_350_60_n_52, sub_350_60_n_54, sub_350_60_n_55,
     sub_350_60_n_56, sub_380_59_n_0, sub_380_59_n_1, sub_380_59_n_2,
     sub_380_59_n_3, sub_380_59_n_4, sub_380_59_n_5, sub_380_59_n_6,
     sub_380_59_n_7, sub_380_59_n_8, sub_380_59_n_10, sub_380_59_n_11,
     sub_380_59_n_12, sub_380_59_n_13, sub_380_59_n_14, sub_380_59_n_15,
     sub_380_59_n_16, sub_380_59_n_17, sub_380_59_n_18, sub_380_59_n_19,
     sub_380_59_n_20, sub_380_59_n_21, sub_380_59_n_22, sub_380_59_n_23,
     sub_380_59_n_24, sub_380_59_n_25, sub_380_59_n_26, sub_380_59_n_27,
     sub_380_59_n_28, sub_380_59_n_29, sub_380_59_n_30, sub_380_59_n_31,
     sub_380_59_n_32, sub_380_59_n_33, sub_380_59_n_34, sub_380_59_n_36,
     sub_380_59_n_37, sub_380_59_n_38, sub_380_59_n_39, sub_380_59_n_40,
     sub_380_59_n_41, sub_380_59_n_42, sub_380_59_n_43, sub_380_59_n_44,
     sub_380_59_n_45, sub_380_59_n_46, sub_380_59_n_47, sub_380_59_n_48,
     sub_380_59_n_49, sub_380_59_n_50, sub_380_59_n_51, sub_380_59_n_52,
     sub_380_59_n_53, sub_380_59_n_54, sub_380_59_n_55, sub_380_59_n_57,
     sub_380_59_n_58, sub_380_59_n_59, sub_380_59_n_61, sub_380_59_n_62,
     sub_380_59_n_63, sub_410_58_n_0, sub_410_58_n_1, sub_410_58_n_2,
     sub_410_58_n_3, sub_410_58_n_4, sub_410_58_n_5, sub_410_58_n_6,
     sub_410_58_n_7, sub_410_58_n_8, sub_410_58_n_9, sub_410_58_n_10,
     sub_410_58_n_11, sub_410_58_n_12, sub_410_58_n_13, sub_410_58_n_14,
     sub_410_58_n_16, sub_410_58_n_17, sub_410_58_n_18, sub_410_58_n_19,
     sub_410_58_n_20, sub_410_58_n_21, sub_410_58_n_22, sub_410_58_n_23,
     sub_410_58_n_24, sub_410_58_n_25, sub_410_58_n_26, sub_410_58_n_27,
     sub_410_58_n_28, sub_410_58_n_29, sub_410_58_n_30, sub_410_58_n_31,
     sub_410_58_n_32, sub_410_58_n_33, sub_410_58_n_34, sub_410_58_n_35,
     sub_410_58_n_36, sub_410_58_n_37, sub_410_58_n_38, sub_410_58_n_39,
     sub_410_58_n_40, sub_410_58_n_41, sub_410_58_n_42, sub_410_58_n_44,
     sub_410_58_n_45, sub_410_58_n_46, sub_410_58_n_47, sub_410_58_n_48,
     sub_410_58_n_49, sub_410_58_n_50, sub_410_58_n_51, sub_410_58_n_52,
     sub_410_58_n_53, sub_410_58_n_54, sub_410_58_n_55, sub_410_58_n_56,
     sub_410_58_n_57, sub_410_58_n_59, sub_410_58_n_60, sub_410_58_n_61,
     sub_410_58_n_62, sub_410_58_n_64, sub_410_58_n_65, sub_410_58_n_67,
     sub_410_58_n_69, sub_440_57_n_0, sub_440_57_n_1, sub_440_57_n_2,
     sub_440_57_n_3, sub_440_57_n_4, sub_440_57_n_5, sub_440_57_n_6,
     sub_440_57_n_7, sub_440_57_n_8, sub_440_57_n_9, sub_440_57_n_10,
     sub_440_57_n_11, sub_440_57_n_12, sub_440_57_n_14, sub_440_57_n_15,
     sub_440_57_n_16, sub_440_57_n_17, sub_440_57_n_18, sub_440_57_n_19,
     sub_440_57_n_20, sub_440_57_n_21, sub_440_57_n_22, sub_440_57_n_23,
     sub_440_57_n_24, sub_440_57_n_25, sub_440_57_n_26, sub_440_57_n_27,
     sub_440_57_n_28, sub_440_57_n_29, sub_440_57_n_30, sub_440_57_n_31,
     sub_440_57_n_32, sub_440_57_n_33, sub_440_57_n_34, sub_440_57_n_35,
     sub_440_57_n_36, sub_440_57_n_37, sub_440_57_n_38, sub_440_57_n_39,
     sub_440_57_n_40, sub_440_57_n_41, sub_440_57_n_43, sub_440_57_n_44,
     sub_440_57_n_45, sub_440_57_n_46, sub_440_57_n_47, sub_440_57_n_48,
     sub_440_57_n_49, sub_440_57_n_50, sub_440_57_n_51, sub_440_57_n_52,
     sub_440_57_n_53, sub_440_57_n_54, sub_440_57_n_55, sub_440_57_n_56,
     sub_440_57_n_57, sub_440_57_n_58, sub_440_57_n_59, sub_440_57_n_60,
     sub_440_57_n_61, sub_440_57_n_62, sub_440_57_n_63, sub_440_57_n_64,
     sub_440_57_n_66, sub_440_57_n_67, sub_440_57_n_68, sub_440_57_n_69,
     sub_440_57_n_70, sub_440_57_n_71, sub_440_57_n_72, sub_440_57_n_73,
     sub_440_57_n_74, sub_440_57_n_76, sub_440_57_n_78, sub_440_57_n_79,
     sub_440_57_n_80, sub_440_57_n_81, sub_470_56_n_0, sub_470_56_n_1,
     sub_470_56_n_2, sub_470_56_n_3, sub_470_56_n_4, sub_470_56_n_5,
     sub_470_56_n_6, sub_470_56_n_7, sub_470_56_n_8, sub_470_56_n_9,
     sub_470_56_n_10, sub_470_56_n_11, sub_470_56_n_12, sub_470_56_n_13,
     sub_470_56_n_15, sub_470_56_n_16, sub_470_56_n_17, sub_470_56_n_18,
     sub_470_56_n_19, sub_470_56_n_20, sub_470_56_n_21, sub_470_56_n_22,
     sub_470_56_n_23, sub_470_56_n_24, sub_470_56_n_25, sub_470_56_n_26,
     sub_470_56_n_27, sub_470_56_n_28, sub_470_56_n_29, sub_470_56_n_31,
     sub_470_56_n_32, sub_470_56_n_33, sub_470_56_n_34, sub_470_56_n_35,
     sub_470_56_n_36, sub_470_56_n_37, sub_470_56_n_38, sub_470_56_n_39,
     sub_470_56_n_40, sub_470_56_n_41, sub_470_56_n_42, sub_470_56_n_43,
     sub_470_56_n_44, sub_470_56_n_46, sub_470_56_n_47, sub_470_56_n_48,
     sub_470_56_n_49, sub_470_56_n_50, sub_470_56_n_51, sub_470_56_n_53,
     sub_470_56_n_54, sub_470_56_n_55, sub_470_56_n_56, sub_470_56_n_59,
     sub_470_56_n_60, sub_470_56_n_61, sub_470_56_n_62, sub_470_56_n_66,
     sub_500_55_n_0, sub_500_55_n_1, sub_500_55_n_2, sub_500_55_n_3,
     sub_500_55_n_4, sub_500_55_n_5, sub_500_55_n_6, sub_500_55_n_7,
     sub_500_55_n_8, sub_500_55_n_9, sub_500_55_n_10, sub_500_55_n_11,
     sub_500_55_n_12, sub_500_55_n_13, sub_500_55_n_14, sub_500_55_n_17,
     sub_500_55_n_18, sub_500_55_n_20, sub_500_55_n_21, sub_500_55_n_22,
     sub_500_55_n_23, sub_500_55_n_24, sub_500_55_n_25, sub_500_55_n_26,
     sub_500_55_n_27, sub_500_55_n_28, sub_500_55_n_29, sub_500_55_n_30,
     sub_500_55_n_31, sub_500_55_n_32, sub_500_55_n_33, sub_500_55_n_34,
     sub_500_55_n_35, sub_500_55_n_36, sub_500_55_n_37, sub_500_55_n_38,
     sub_500_55_n_39, sub_500_55_n_40, sub_500_55_n_41, sub_500_55_n_42,
     sub_500_55_n_43, sub_500_55_n_44, sub_500_55_n_45, sub_500_55_n_47,
     sub_500_55_n_48, sub_500_55_n_49, sub_500_55_n_50, sub_500_55_n_51,
     sub_500_55_n_52, sub_500_55_n_53, sub_500_55_n_54, sub_500_55_n_55,
     sub_500_55_n_56, sub_500_55_n_57, sub_500_55_n_58, sub_500_55_n_59,
     sub_500_55_n_60, sub_500_55_n_61, sub_500_55_n_62, sub_500_55_n_63,
     sub_500_55_n_64, sub_500_55_n_66, sub_500_55_n_67, sub_500_55_n_68,
     sub_500_55_n_69, sub_500_55_n_70, sub_500_55_n_72, sub_500_55_n_73,
     sub_500_55_n_74, sub_500_55_n_75, sub_500_55_n_77, sub_500_55_n_78,
     sub_500_55_n_79, sub_500_55_n_80, sub_500_55_n_81, sub_500_55_n_85,
     sub_530_54_n_0, sub_530_54_n_1, sub_530_54_n_2, sub_530_54_n_3,
     sub_530_54_n_4, sub_530_54_n_5, sub_530_54_n_6, sub_530_54_n_7,
     sub_530_54_n_8, sub_530_54_n_9, sub_530_54_n_10, sub_530_54_n_11,
     sub_530_54_n_12, sub_530_54_n_13, sub_530_54_n_14, sub_530_54_n_16,
     sub_530_54_n_17, sub_530_54_n_18, sub_530_54_n_19, sub_530_54_n_20,
     sub_530_54_n_21, sub_530_54_n_23, sub_530_54_n_24, sub_530_54_n_25,
     sub_530_54_n_26, sub_530_54_n_27, sub_530_54_n_28, sub_530_54_n_29,
     sub_530_54_n_30, sub_530_54_n_31, sub_530_54_n_32, sub_530_54_n_33,
     sub_530_54_n_34, sub_530_54_n_35, sub_530_54_n_36, sub_530_54_n_37,
     sub_530_54_n_38, sub_530_54_n_39, sub_530_54_n_40, sub_530_54_n_41,
     sub_530_54_n_42, sub_530_54_n_43, sub_530_54_n_44, sub_530_54_n_45,
     sub_530_54_n_46, sub_530_54_n_48, sub_530_54_n_49, sub_530_54_n_50,
     sub_530_54_n_51, sub_530_54_n_52, sub_530_54_n_53, sub_530_54_n_54,
     sub_530_54_n_55, sub_530_54_n_56, sub_530_54_n_57, sub_530_54_n_58,
     sub_530_54_n_59, sub_530_54_n_60, sub_530_54_n_61, sub_530_54_n_62,
     sub_530_54_n_63, sub_530_54_n_64, sub_530_54_n_65, sub_530_54_n_67,
     sub_530_54_n_68, sub_530_54_n_69, sub_530_54_n_70, sub_530_54_n_71,
     sub_530_54_n_72, sub_530_54_n_73, sub_530_54_n_74, sub_530_54_n_76,
     sub_530_54_n_77, sub_530_54_n_78, sub_530_54_n_79, sub_530_54_n_81,
     sub_530_54_n_82, sub_530_54_n_87, sub_530_54_n_88, sub_530_54_n_89,
     sub_560_53_n_0, sub_560_53_n_1, sub_560_53_n_2, sub_560_53_n_3,
     sub_560_53_n_4, sub_560_53_n_5, sub_560_53_n_6, sub_560_53_n_7,
     sub_560_53_n_8, sub_560_53_n_9, sub_560_53_n_10, sub_560_53_n_11,
     sub_560_53_n_12, sub_560_53_n_13, sub_560_53_n_14, sub_560_53_n_15,
     sub_560_53_n_16, sub_560_53_n_17, sub_560_53_n_18, sub_560_53_n_19,
     sub_560_53_n_20, sub_560_53_n_21, sub_560_53_n_23, sub_560_53_n_24,
     sub_560_53_n_25, sub_560_53_n_26, sub_560_53_n_27, sub_560_53_n_28,
     sub_560_53_n_29, sub_560_53_n_30, sub_560_53_n_31, sub_560_53_n_32,
     sub_560_53_n_33, sub_560_53_n_34, sub_560_53_n_35, sub_560_53_n_36,
     sub_560_53_n_37, sub_560_53_n_38, sub_560_53_n_39, sub_560_53_n_40,
     sub_560_53_n_41, sub_560_53_n_42, sub_560_53_n_43, sub_560_53_n_44,
     sub_560_53_n_45, sub_560_53_n_46, sub_560_53_n_48, sub_560_53_n_49,
     sub_560_53_n_50, sub_560_53_n_51, sub_560_53_n_52, sub_560_53_n_53,
     sub_560_53_n_54, sub_560_53_n_55, sub_560_53_n_56, sub_560_53_n_57,
     sub_560_53_n_58, sub_560_53_n_59, sub_560_53_n_60, sub_560_53_n_61,
     sub_560_53_n_62, sub_560_53_n_63, sub_560_53_n_64, sub_560_53_n_65,
     sub_560_53_n_66, sub_560_53_n_67, sub_560_53_n_68, sub_560_53_n_69,
     sub_560_53_n_70, sub_560_53_n_71, sub_560_53_n_72, sub_560_53_n_73,
     sub_560_53_n_75, sub_560_53_n_76, sub_560_53_n_77, sub_560_53_n_78,
     sub_560_53_n_79, sub_560_53_n_81, sub_560_53_n_82, sub_560_53_n_83,
     sub_560_53_n_84, sub_560_53_n_85, sub_560_53_n_87, sub_560_53_n_88,
     sub_560_53_n_89, sub_560_53_n_91, sub_560_53_n_95, sub_560_53_n_96,
     sub_560_53_n_97, sub_560_53_n_98, sub_560_53_n_103, sub_590_52_n_0,
     sub_590_52_n_1, sub_590_52_n_2, sub_590_52_n_3, sub_590_52_n_4,
     sub_590_52_n_5, sub_590_52_n_6, sub_590_52_n_7, sub_590_52_n_8,
     sub_590_52_n_9, sub_590_52_n_10, sub_590_52_n_11, sub_590_52_n_12,
     sub_590_52_n_13, sub_590_52_n_14, sub_590_52_n_15, sub_590_52_n_16,
     sub_590_52_n_17, sub_590_52_n_20, sub_590_52_n_21, sub_590_52_n_22,
     sub_590_52_n_23, sub_590_52_n_24, sub_590_52_n_25, sub_590_52_n_26,
     sub_590_52_n_28, sub_590_52_n_29, sub_590_52_n_30, sub_590_52_n_31,
     sub_590_52_n_32, sub_590_52_n_33, sub_590_52_n_34, sub_590_52_n_35,
     sub_590_52_n_36, sub_590_52_n_37, sub_590_52_n_38, sub_590_52_n_39,
     sub_590_52_n_40, sub_590_52_n_41, sub_590_52_n_42, sub_590_52_n_43,
     sub_590_52_n_44, sub_590_52_n_45, sub_590_52_n_46, sub_590_52_n_47,
     sub_590_52_n_48, sub_590_52_n_49, sub_590_52_n_50, sub_590_52_n_51,
     sub_590_52_n_52, sub_590_52_n_53, sub_590_52_n_54, sub_590_52_n_55,
     sub_590_52_n_56, sub_590_52_n_57, sub_590_52_n_59, sub_590_52_n_60,
     sub_590_52_n_61, sub_590_52_n_62, sub_590_52_n_63, sub_590_52_n_64,
     sub_590_52_n_65, sub_590_52_n_66, sub_590_52_n_67, sub_590_52_n_68,
     sub_590_52_n_69, sub_590_52_n_70, sub_590_52_n_71, sub_590_52_n_72,
     sub_590_52_n_73, sub_590_52_n_74, sub_590_52_n_75, sub_590_52_n_76,
     sub_590_52_n_77, sub_590_52_n_78, sub_590_52_n_80, sub_590_52_n_81,
     sub_590_52_n_82, sub_590_52_n_83, sub_590_52_n_84, sub_590_52_n_85,
     sub_590_52_n_86, sub_590_52_n_87, sub_590_52_n_89, sub_590_52_n_90,
     sub_590_52_n_92, sub_590_52_n_93, sub_590_52_n_94, sub_590_52_n_95,
     sub_590_52_n_96, sub_590_52_n_97, sub_590_52_n_100, sub_590_52_n_101,
     sub_590_52_n_104, sub_590_52_n_105, sub_620_51_n_0, sub_620_51_n_1,
     sub_620_51_n_2, sub_620_51_n_3, sub_620_51_n_4, sub_620_51_n_5,
     sub_620_51_n_6, sub_620_51_n_7, sub_620_51_n_8, sub_620_51_n_9,
     sub_620_51_n_10, sub_620_51_n_11, sub_620_51_n_12, sub_620_51_n_13,
     sub_620_51_n_14, sub_620_51_n_15, sub_620_51_n_16, sub_620_51_n_17,
     sub_620_51_n_18, sub_620_51_n_19, sub_620_51_n_20, sub_620_51_n_22,
     sub_620_51_n_23, sub_620_51_n_24, sub_620_51_n_25, sub_620_51_n_26,
     sub_620_51_n_27, sub_620_51_n_28, sub_620_51_n_29, sub_620_51_n_30,
     sub_620_51_n_32, sub_620_51_n_33, sub_620_51_n_34, sub_620_51_n_35,
     sub_620_51_n_36, sub_620_51_n_37, sub_620_51_n_38, sub_620_51_n_39,
     sub_620_51_n_40, sub_620_51_n_41, sub_620_51_n_42, sub_620_51_n_43,
     sub_620_51_n_44, sub_620_51_n_45, sub_620_51_n_46, sub_620_51_n_47,
     sub_620_51_n_48, sub_620_51_n_49, sub_620_51_n_50, sub_620_51_n_51,
     sub_620_51_n_52, sub_620_51_n_53, sub_620_51_n_54, sub_620_51_n_55,
     sub_620_51_n_56, sub_620_51_n_57, sub_620_51_n_58, sub_620_51_n_60,
     sub_620_51_n_61, sub_620_51_n_62, sub_620_51_n_63, sub_620_51_n_64,
     sub_620_51_n_65, sub_620_51_n_66, sub_620_51_n_67, sub_620_51_n_68,
     sub_620_51_n_69, sub_620_51_n_70, sub_620_51_n_71, sub_620_51_n_72,
     sub_620_51_n_73, sub_620_51_n_74, sub_620_51_n_75, sub_620_51_n_76,
     sub_620_51_n_77, sub_620_51_n_78, sub_620_51_n_79, sub_620_51_n_80,
     sub_620_51_n_81, sub_620_51_n_82, sub_620_51_n_83, sub_620_51_n_84,
     sub_620_51_n_85, sub_620_51_n_86, sub_620_51_n_88, sub_620_51_n_89,
     sub_620_51_n_90, sub_620_51_n_91, sub_620_51_n_92, sub_620_51_n_93,
     sub_620_51_n_94, sub_620_51_n_96, sub_620_51_n_97, sub_620_51_n_98,
     sub_620_51_n_100, sub_620_51_n_101, sub_620_51_n_103, sub_620_51_n_106,
     sub_620_51_n_107, sub_620_51_n_108, sub_620_51_n_111, sub_620_51_n_115,
     sub_650_50_n_0, sub_650_50_n_1, sub_650_50_n_2, sub_650_50_n_3,
     sub_650_50_n_4, sub_650_50_n_5, sub_650_50_n_6, sub_650_50_n_7,
     sub_650_50_n_8, sub_650_50_n_9, sub_650_50_n_10, sub_650_50_n_11,
     sub_650_50_n_12, sub_650_50_n_13, sub_650_50_n_14, sub_650_50_n_15,
     sub_650_50_n_16, sub_650_50_n_17, sub_650_50_n_18, sub_650_50_n_19,
     sub_650_50_n_20, sub_650_50_n_21, sub_650_50_n_22, sub_650_50_n_23,
     sub_650_50_n_24, sub_650_50_n_26, sub_650_50_n_27, sub_650_50_n_28,
     sub_650_50_n_29, sub_650_50_n_30, sub_650_50_n_31, sub_650_50_n_32,
     sub_650_50_n_33, sub_650_50_n_34, sub_650_50_n_35, sub_650_50_n_36,
     sub_650_50_n_37, sub_650_50_n_39, sub_650_50_n_40, sub_650_50_n_41,
     sub_650_50_n_42, sub_650_50_n_43, sub_650_50_n_44, sub_650_50_n_45,
     sub_650_50_n_46, sub_650_50_n_47, sub_650_50_n_48, sub_650_50_n_49,
     sub_650_50_n_50, sub_650_50_n_51, sub_650_50_n_52, sub_650_50_n_53,
     sub_650_50_n_54, sub_650_50_n_55, sub_650_50_n_56, sub_650_50_n_57,
     sub_650_50_n_58, sub_650_50_n_59, sub_650_50_n_60, sub_650_50_n_61,
     sub_650_50_n_62, sub_650_50_n_64, sub_650_50_n_65, sub_650_50_n_66,
     sub_650_50_n_67, sub_650_50_n_68, sub_650_50_n_69, sub_650_50_n_70,
     sub_650_50_n_71, sub_650_50_n_72, sub_650_50_n_73, sub_650_50_n_74,
     sub_650_50_n_75, sub_650_50_n_76, sub_650_50_n_77, sub_650_50_n_78,
     sub_650_50_n_79, sub_650_50_n_80, sub_650_50_n_81, sub_650_50_n_82,
     sub_650_50_n_83, sub_650_50_n_84, sub_650_50_n_85, sub_650_50_n_86,
     sub_650_50_n_87, sub_650_50_n_88, sub_650_50_n_89, sub_650_50_n_90,
     sub_650_50_n_91, sub_650_50_n_92, sub_650_50_n_93, sub_650_50_n_94,
     sub_650_50_n_95, sub_650_50_n_97, sub_650_50_n_98, sub_650_50_n_99,
     sub_650_50_n_100, sub_650_50_n_101, sub_650_50_n_102, sub_650_50_n_103,
     sub_650_50_n_104, sub_650_50_n_106, sub_650_50_n_107, sub_650_50_n_108,
     sub_650_50_n_110, sub_650_50_n_111, sub_650_50_n_112, sub_650_50_n_116,
     sub_650_50_n_117, sub_650_50_n_118, sub_650_50_n_119, sub_650_50_n_120,
     sub_650_50_n_126, sub_680_49_n_0, sub_680_49_n_1, sub_680_49_n_2,
     sub_680_49_n_3, sub_680_49_n_4, sub_680_49_n_5, sub_680_49_n_6,
     sub_680_49_n_7, sub_680_49_n_8, sub_680_49_n_9, sub_680_49_n_10,
     sub_680_49_n_11, sub_680_49_n_12, sub_680_49_n_13, sub_680_49_n_14,
     sub_680_49_n_16, sub_680_49_n_17, sub_680_49_n_18, sub_680_49_n_19,
     sub_680_49_n_20, sub_680_49_n_21, sub_680_49_n_22, sub_680_49_n_23,
     sub_680_49_n_24, sub_680_49_n_25, sub_680_49_n_27, sub_680_49_n_28,
     sub_680_49_n_29, sub_680_49_n_30, sub_680_49_n_31, sub_680_49_n_32,
     sub_680_49_n_33, sub_680_49_n_34, sub_680_49_n_35, sub_680_49_n_36,
     sub_680_49_n_37, sub_680_49_n_38, sub_680_49_n_39, sub_680_49_n_40,
     sub_680_49_n_41, sub_680_49_n_42, sub_680_49_n_43, sub_680_49_n_44,
     sub_680_49_n_45, sub_680_49_n_46, sub_680_49_n_47, sub_680_49_n_48,
     sub_680_49_n_49, sub_680_49_n_50, sub_680_49_n_51, sub_680_49_n_52,
     sub_680_49_n_53, sub_680_49_n_54, sub_680_49_n_55, sub_680_49_n_56,
     sub_680_49_n_57, sub_680_49_n_58, sub_680_49_n_59, sub_680_49_n_60,
     sub_680_49_n_61, sub_680_49_n_62, sub_680_49_n_63, sub_680_49_n_64,
     sub_680_49_n_65, sub_680_49_n_67, sub_680_49_n_68, sub_680_49_n_69,
     sub_680_49_n_70, sub_680_49_n_71, sub_680_49_n_72, sub_680_49_n_73,
     sub_680_49_n_74, sub_680_49_n_75, sub_680_49_n_76, sub_680_49_n_77,
     sub_680_49_n_78, sub_680_49_n_79, sub_680_49_n_80, sub_680_49_n_81,
     sub_680_49_n_82, sub_680_49_n_83, sub_680_49_n_84, sub_680_49_n_85,
     sub_680_49_n_86, sub_680_49_n_87, sub_680_49_n_88, sub_680_49_n_89,
     sub_680_49_n_90, sub_680_49_n_91, sub_680_49_n_92, sub_680_49_n_93,
     sub_680_49_n_94, sub_680_49_n_95, sub_680_49_n_96, sub_680_49_n_97,
     sub_680_49_n_98, sub_680_49_n_99, sub_680_49_n_100, sub_680_49_n_101,
     sub_680_49_n_102, sub_680_49_n_103, sub_680_49_n_104, sub_680_49_n_105,
     sub_680_49_n_106, sub_680_49_n_107, sub_680_49_n_108, sub_680_49_n_110,
     sub_680_49_n_111, sub_680_49_n_112, sub_680_49_n_113, sub_680_49_n_115,
     sub_680_49_n_116, sub_680_49_n_117, sub_680_49_n_118, sub_680_49_n_119,
     sub_680_49_n_120, sub_680_49_n_121, sub_680_49_n_123, sub_680_49_n_124,
     sub_680_49_n_125, sub_680_49_n_126, sub_680_49_n_127, sub_680_49_n_128,
     sub_680_49_n_132, sub_680_49_n_133, sub_680_49_n_134, sub_680_49_n_135,
     sub_680_49_n_136, sub_680_49_n_143, sub_680_49_n_144, sub_710_48_n_0,
     sub_710_48_n_1, sub_710_48_n_2, sub_710_48_n_3, sub_710_48_n_4,
     sub_710_48_n_5, sub_710_48_n_6, sub_710_48_n_7, sub_710_48_n_8,
     sub_710_48_n_9, sub_710_48_n_10, sub_710_48_n_11, sub_710_48_n_12,
     sub_710_48_n_13, sub_710_48_n_14, sub_710_48_n_15, sub_710_48_n_16,
     sub_710_48_n_17, sub_710_48_n_18, sub_710_48_n_19, sub_710_48_n_20,
     sub_710_48_n_21, sub_710_48_n_22, sub_710_48_n_23, sub_710_48_n_24,
     sub_710_48_n_25, sub_710_48_n_26, sub_710_48_n_27, sub_710_48_n_28,
     sub_710_48_n_29, sub_710_48_n_30, sub_710_48_n_31, sub_710_48_n_32,
     sub_710_48_n_33, sub_710_48_n_34, sub_710_48_n_36, sub_710_48_n_37,
     sub_710_48_n_38, sub_710_48_n_39, sub_710_48_n_40, sub_710_48_n_41,
     sub_710_48_n_42, sub_710_48_n_43, sub_710_48_n_44, sub_710_48_n_45,
     sub_710_48_n_46, sub_710_48_n_47, sub_710_48_n_48, sub_710_48_n_49,
     sub_710_48_n_50, sub_710_48_n_51, sub_710_48_n_52, sub_710_48_n_53,
     sub_710_48_n_54, sub_710_48_n_55, sub_710_48_n_56, sub_710_48_n_57,
     sub_710_48_n_58, sub_710_48_n_59, sub_710_48_n_60, sub_710_48_n_61,
     sub_710_48_n_62, sub_710_48_n_63, sub_710_48_n_64, sub_710_48_n_65,
     sub_710_48_n_66, sub_710_48_n_67, sub_710_48_n_69, sub_710_48_n_70,
     sub_710_48_n_71, sub_710_48_n_72, sub_710_48_n_73, sub_710_48_n_74,
     sub_710_48_n_75, sub_710_48_n_76, sub_710_48_n_77, sub_710_48_n_78,
     sub_710_48_n_79, sub_710_48_n_80, sub_710_48_n_81, sub_710_48_n_82,
     sub_710_48_n_83, sub_710_48_n_84, sub_710_48_n_85, sub_710_48_n_86,
     sub_710_48_n_87, sub_710_48_n_88, sub_710_48_n_89, sub_710_48_n_90,
     sub_710_48_n_91, sub_710_48_n_92, sub_710_48_n_93, sub_710_48_n_94,
     sub_710_48_n_95, sub_710_48_n_96, sub_710_48_n_97, sub_710_48_n_98,
     sub_710_48_n_99, sub_710_48_n_100, sub_710_48_n_101, sub_710_48_n_102,
     sub_710_48_n_103, sub_710_48_n_104, sub_710_48_n_105, sub_710_48_n_106,
     sub_710_48_n_107, sub_710_48_n_108, sub_710_48_n_109, sub_710_48_n_110,
     sub_710_48_n_111, sub_710_48_n_113, sub_710_48_n_114, sub_710_48_n_115,
     sub_710_48_n_116, sub_710_48_n_117, sub_710_48_n_119, sub_710_48_n_120,
     sub_710_48_n_121, sub_710_48_n_122, sub_710_48_n_123, sub_710_48_n_126,
     sub_710_48_n_127, sub_710_48_n_128, sub_710_48_n_129, sub_710_48_n_130,
     sub_710_48_n_132, sub_710_48_n_133, sub_710_48_n_134, sub_710_48_n_137,
     sub_710_48_n_138, sub_710_48_n_139, sub_710_48_n_140, sub_710_48_n_141,
     sub_710_48_n_142, sub_710_48_n_146, sub_710_48_n_147, sub_710_48_n_148,
     sub_710_48_n_149, sub_710_48_n_153, sub_740_47_n_0, sub_740_47_n_1,
     sub_740_47_n_2, sub_740_47_n_3, sub_740_47_n_4, sub_740_47_n_5,
     sub_740_47_n_6, sub_740_47_n_7, sub_740_47_n_8, sub_740_47_n_9,
     sub_740_47_n_10, sub_740_47_n_11, sub_740_47_n_12, sub_740_47_n_13,
     sub_740_47_n_14, sub_740_47_n_15, sub_740_47_n_16, sub_740_47_n_17,
     sub_740_47_n_18, sub_740_47_n_19, sub_740_47_n_20, sub_740_47_n_21,
     sub_740_47_n_22, sub_740_47_n_23, sub_740_47_n_24, sub_740_47_n_25,
     sub_740_47_n_26, sub_740_47_n_27, sub_740_47_n_28, sub_740_47_n_29,
     sub_740_47_n_30, sub_740_47_n_31, sub_740_47_n_32, sub_740_47_n_33,
     sub_740_47_n_34, sub_740_47_n_35, sub_740_47_n_36, sub_740_47_n_37,
     sub_740_47_n_38, sub_740_47_n_39, sub_740_47_n_40, sub_740_47_n_41,
     sub_740_47_n_42, sub_740_47_n_43, sub_740_47_n_45, sub_740_47_n_46,
     sub_740_47_n_47, sub_740_47_n_48, sub_740_47_n_49, sub_740_47_n_50,
     sub_740_47_n_51, sub_740_47_n_52, sub_740_47_n_53, sub_740_47_n_54,
     sub_740_47_n_55, sub_740_47_n_56, sub_740_47_n_57, sub_740_47_n_58,
     sub_740_47_n_59, sub_740_47_n_60, sub_740_47_n_61, sub_740_47_n_62,
     sub_740_47_n_63, sub_740_47_n_64, sub_740_47_n_65, sub_740_47_n_66,
     sub_740_47_n_67, sub_740_47_n_68, sub_740_47_n_69, sub_740_47_n_70,
     sub_740_47_n_71, sub_740_47_n_72, sub_740_47_n_74, sub_740_47_n_75,
     sub_740_47_n_76, sub_740_47_n_77, sub_740_47_n_78, sub_740_47_n_79,
     sub_740_47_n_80, sub_740_47_n_81, sub_740_47_n_82, sub_740_47_n_83,
     sub_740_47_n_84, sub_740_47_n_85, sub_740_47_n_86, sub_740_47_n_87,
     sub_740_47_n_88, sub_740_47_n_89, sub_740_47_n_90, sub_740_47_n_91,
     sub_740_47_n_92, sub_740_47_n_93, sub_740_47_n_94, sub_740_47_n_95,
     sub_740_47_n_96, sub_740_47_n_97, sub_740_47_n_98, sub_740_47_n_99,
     sub_740_47_n_100, sub_740_47_n_101, sub_740_47_n_102, sub_740_47_n_104,
     sub_740_47_n_105, sub_740_47_n_106, sub_740_47_n_108, sub_740_47_n_109,
     sub_740_47_n_110, sub_740_47_n_113, sub_740_47_n_114, sub_740_47_n_115,
     sub_740_47_n_116, sub_740_47_n_117, sub_740_47_n_118, sub_740_47_n_122,
     sub_740_47_n_123, sub_740_47_n_124, sub_740_47_n_125, sub_740_47_n_126,
     sub_740_47_n_127, sub_740_47_n_133, sub_740_47_n_134, sub_740_47_n_135,
     sub_740_47_n_136, sub_740_47_n_138, sub_740_47_n_143, sub_770_46_n_0,
     sub_770_46_n_1, sub_770_46_n_2, sub_770_46_n_3, sub_770_46_n_4,
     sub_770_46_n_5, sub_770_46_n_6, sub_770_46_n_7, sub_770_46_n_8,
     sub_770_46_n_9, sub_770_46_n_10, sub_770_46_n_11, sub_770_46_n_12,
     sub_770_46_n_13, sub_770_46_n_14, sub_770_46_n_15, sub_770_46_n_16,
     sub_770_46_n_17, sub_770_46_n_18, sub_770_46_n_19, sub_770_46_n_20,
     sub_770_46_n_21, sub_770_46_n_22, sub_770_46_n_23, sub_770_46_n_24,
     sub_770_46_n_26, sub_770_46_n_28, sub_770_46_n_29, sub_770_46_n_31,
     sub_770_46_n_32, sub_770_46_n_33, sub_770_46_n_34, sub_770_46_n_35,
     sub_770_46_n_36, sub_770_46_n_37, sub_770_46_n_38, sub_770_46_n_39,
     sub_770_46_n_40, sub_770_46_n_42, sub_770_46_n_43, sub_770_46_n_44,
     sub_770_46_n_45, sub_770_46_n_46, sub_770_46_n_47, sub_770_46_n_48,
     sub_770_46_n_49, sub_770_46_n_50, sub_770_46_n_51, sub_770_46_n_52,
     sub_770_46_n_53, sub_770_46_n_54, sub_770_46_n_55, sub_770_46_n_56,
     sub_770_46_n_57, sub_770_46_n_58, sub_770_46_n_59, sub_770_46_n_60,
     sub_770_46_n_61, sub_770_46_n_62, sub_770_46_n_63, sub_770_46_n_64,
     sub_770_46_n_65, sub_770_46_n_66, sub_770_46_n_67, sub_770_46_n_68,
     sub_770_46_n_69, sub_770_46_n_70, sub_770_46_n_72, sub_770_46_n_73,
     sub_770_46_n_74, sub_770_46_n_75, sub_770_46_n_76, sub_770_46_n_77,
     sub_770_46_n_78, sub_770_46_n_79, sub_770_46_n_80, sub_770_46_n_81,
     sub_770_46_n_82, sub_770_46_n_83, sub_770_46_n_84, sub_770_46_n_85,
     sub_770_46_n_86, sub_770_46_n_87, sub_770_46_n_88, sub_770_46_n_89,
     sub_770_46_n_90, sub_770_46_n_91, sub_770_46_n_92, sub_770_46_n_93,
     sub_770_46_n_94, sub_770_46_n_95, sub_770_46_n_96, sub_770_46_n_97,
     sub_770_46_n_98, sub_770_46_n_99, sub_770_46_n_100, sub_770_46_n_101,
     sub_770_46_n_102, sub_770_46_n_103, sub_770_46_n_104, sub_770_46_n_105,
     sub_770_46_n_106, sub_770_46_n_107, sub_770_46_n_108, sub_770_46_n_109,
     sub_770_46_n_110, sub_770_46_n_111, sub_770_46_n_112, sub_770_46_n_114,
     sub_770_46_n_115, sub_770_46_n_116, sub_770_46_n_118, sub_770_46_n_119,
     sub_770_46_n_120, sub_770_46_n_123, sub_770_46_n_124, sub_770_46_n_125,
     sub_770_46_n_126, sub_770_46_n_127, sub_770_46_n_129, sub_770_46_n_130,
     sub_770_46_n_131, sub_770_46_n_132, sub_770_46_n_133, sub_770_46_n_134,
     sub_770_46_n_135, sub_770_46_n_136, sub_770_46_n_141, sub_770_46_n_142,
     sub_770_46_n_143, sub_770_46_n_144, sub_770_46_n_145, sub_800_45_n_0,
     sub_800_45_n_1, sub_800_45_n_2, sub_800_45_n_3, sub_800_45_n_4,
     sub_800_45_n_5, sub_800_45_n_6, sub_800_45_n_7, sub_800_45_n_8,
     sub_800_45_n_9, sub_800_45_n_10, sub_800_45_n_11, sub_800_45_n_12,
     sub_800_45_n_13, sub_800_45_n_14, sub_800_45_n_15, sub_800_45_n_16,
     sub_800_45_n_17, sub_800_45_n_18, sub_800_45_n_19, sub_800_45_n_20,
     sub_800_45_n_21, sub_800_45_n_22, sub_800_45_n_23, sub_800_45_n_24,
     sub_800_45_n_25, sub_800_45_n_26, sub_800_45_n_27, sub_800_45_n_28,
     sub_800_45_n_29, sub_800_45_n_30, sub_800_45_n_31, sub_800_45_n_32,
     sub_800_45_n_34, sub_800_45_n_35, sub_800_45_n_36, sub_800_45_n_37,
     sub_800_45_n_38, sub_800_45_n_39, sub_800_45_n_40, sub_800_45_n_41,
     sub_800_45_n_42, sub_800_45_n_43, sub_800_45_n_44, sub_800_45_n_45,
     sub_800_45_n_46, sub_800_45_n_47, sub_800_45_n_48, sub_800_45_n_49,
     sub_800_45_n_50, sub_800_45_n_51, sub_800_45_n_52, sub_800_45_n_53,
     sub_800_45_n_54, sub_800_45_n_55, sub_800_45_n_56, sub_800_45_n_57,
     sub_800_45_n_58, sub_800_45_n_59, sub_800_45_n_60, sub_800_45_n_61,
     sub_800_45_n_62, sub_800_45_n_63, sub_800_45_n_64, sub_800_45_n_65,
     sub_800_45_n_66, sub_800_45_n_67, sub_800_45_n_68, sub_800_45_n_69,
     sub_800_45_n_70, sub_800_45_n_71, sub_800_45_n_73, sub_800_45_n_74,
     sub_800_45_n_75, sub_800_45_n_76, sub_800_45_n_77, sub_800_45_n_78,
     sub_800_45_n_79, sub_800_45_n_80, sub_800_45_n_81, sub_800_45_n_82,
     sub_800_45_n_83, sub_800_45_n_84, sub_800_45_n_85, sub_800_45_n_86,
     sub_800_45_n_87, sub_800_45_n_88, sub_800_45_n_89, sub_800_45_n_90,
     sub_800_45_n_91, sub_800_45_n_92, sub_800_45_n_93, sub_800_45_n_94,
     sub_800_45_n_95, sub_800_45_n_96, sub_800_45_n_97, sub_800_45_n_98,
     sub_800_45_n_99, sub_800_45_n_100, sub_800_45_n_101, sub_800_45_n_102,
     sub_800_45_n_103, sub_800_45_n_104, sub_800_45_n_105, sub_800_45_n_106,
     sub_800_45_n_107, sub_800_45_n_108, sub_800_45_n_109, sub_800_45_n_111,
     sub_800_45_n_112, sub_800_45_n_113, sub_800_45_n_114, sub_800_45_n_115,
     sub_800_45_n_116, sub_800_45_n_117, sub_800_45_n_118, sub_800_45_n_119,
     sub_800_45_n_120, sub_800_45_n_121, sub_800_45_n_123, sub_800_45_n_124,
     sub_800_45_n_125, sub_800_45_n_128, sub_800_45_n_129, sub_800_45_n_130,
     sub_800_45_n_131, sub_800_45_n_132, sub_800_45_n_133, sub_800_45_n_134,
     sub_800_45_n_138, sub_800_45_n_139, sub_800_45_n_140, sub_800_45_n_141,
     sub_800_45_n_142, sub_800_45_n_143, sub_800_45_n_144, sub_800_45_n_145,
     sub_800_45_n_146, sub_800_45_n_147, sub_800_45_n_153, sub_800_45_n_155,
     sub_800_45_n_156, sub_800_45_n_157, sub_800_45_n_158, sub_800_45_n_159,
     sub_800_45_n_160, sub_800_45_n_161, sub_800_45_n_167, sub_800_45_n_168,
     sub_800_45_n_169, sub_830_44_n_0, sub_830_44_n_1, sub_830_44_n_2,
     sub_830_44_n_3, sub_830_44_n_4, sub_830_44_n_5, sub_830_44_n_6,
     sub_830_44_n_7, sub_830_44_n_8, sub_830_44_n_9, sub_830_44_n_10,
     sub_830_44_n_11, sub_830_44_n_12, sub_830_44_n_13, sub_830_44_n_14,
     sub_830_44_n_15, sub_830_44_n_16, sub_830_44_n_17, sub_830_44_n_18,
     sub_830_44_n_19, sub_830_44_n_20, sub_830_44_n_21, sub_830_44_n_22,
     sub_830_44_n_23, sub_830_44_n_24, sub_830_44_n_25, sub_830_44_n_26,
     sub_830_44_n_27, sub_830_44_n_28, sub_830_44_n_29, sub_830_44_n_30,
     sub_830_44_n_31, sub_830_44_n_33, sub_830_44_n_34, sub_830_44_n_35,
     sub_830_44_n_36, sub_830_44_n_37, sub_830_44_n_38, sub_830_44_n_39,
     sub_830_44_n_40, sub_830_44_n_41, sub_830_44_n_42, sub_830_44_n_43,
     sub_830_44_n_44, sub_830_44_n_45, sub_830_44_n_46, sub_830_44_n_47,
     sub_830_44_n_49, sub_830_44_n_50, sub_830_44_n_51, sub_830_44_n_52,
     sub_830_44_n_53, sub_830_44_n_54, sub_830_44_n_55, sub_830_44_n_56,
     sub_830_44_n_57, sub_830_44_n_58, sub_830_44_n_59, sub_830_44_n_60,
     sub_830_44_n_61, sub_830_44_n_62, sub_830_44_n_63, sub_830_44_n_64,
     sub_830_44_n_65, sub_830_44_n_66, sub_830_44_n_67, sub_830_44_n_68,
     sub_830_44_n_69, sub_830_44_n_70, sub_830_44_n_71, sub_830_44_n_72,
     sub_830_44_n_73, sub_830_44_n_74, sub_830_44_n_75, sub_830_44_n_76,
     sub_830_44_n_77, sub_830_44_n_78, sub_830_44_n_79, sub_830_44_n_80,
     sub_830_44_n_81, sub_830_44_n_82, sub_830_44_n_83, sub_830_44_n_84,
     sub_830_44_n_85, sub_830_44_n_86, sub_830_44_n_87, sub_830_44_n_88,
     sub_830_44_n_89, sub_830_44_n_90, sub_830_44_n_92, sub_830_44_n_93,
     sub_830_44_n_94, sub_830_44_n_95, sub_830_44_n_96, sub_830_44_n_97,
     sub_830_44_n_98, sub_830_44_n_99, sub_830_44_n_100, sub_830_44_n_101,
     sub_830_44_n_102, sub_830_44_n_103, sub_830_44_n_104, sub_830_44_n_105,
     sub_830_44_n_106, sub_830_44_n_107, sub_830_44_n_108, sub_830_44_n_109,
     sub_830_44_n_110, sub_830_44_n_111, sub_830_44_n_112, sub_830_44_n_113,
     sub_830_44_n_114, sub_830_44_n_115, sub_830_44_n_116, sub_830_44_n_117,
     sub_830_44_n_118, sub_830_44_n_119, sub_830_44_n_120, sub_830_44_n_121,
     sub_830_44_n_122, sub_830_44_n_123, sub_830_44_n_124, sub_830_44_n_125,
     sub_830_44_n_126, sub_830_44_n_127, sub_830_44_n_128, sub_830_44_n_129,
     sub_830_44_n_130, sub_830_44_n_131, sub_830_44_n_132, sub_830_44_n_133,
     sub_830_44_n_134, sub_830_44_n_135, sub_830_44_n_136, sub_830_44_n_137,
     sub_830_44_n_138, sub_830_44_n_140, sub_830_44_n_141, sub_830_44_n_142,
     sub_830_44_n_144, sub_830_44_n_145, sub_830_44_n_146, sub_830_44_n_147,
     sub_830_44_n_150, sub_830_44_n_151, sub_830_44_n_152, sub_830_44_n_153,
     sub_830_44_n_154, sub_830_44_n_157, sub_830_44_n_158, sub_830_44_n_159,
     sub_830_44_n_160, sub_830_44_n_161, sub_830_44_n_162, sub_830_44_n_163,
     sub_830_44_n_164, sub_830_44_n_165, sub_830_44_n_171, sub_830_44_n_172,
     sub_830_44_n_173, sub_830_44_n_174, sub_830_44_n_182, sub_860_43_n_0,
     sub_860_43_n_1, sub_860_43_n_2, sub_860_43_n_3, sub_860_43_n_4,
     sub_860_43_n_5, sub_860_43_n_6, sub_860_43_n_7, sub_860_43_n_8,
     sub_860_43_n_9, sub_860_43_n_10, sub_860_43_n_11, sub_860_43_n_12,
     sub_860_43_n_13, sub_860_43_n_14, sub_860_43_n_15, sub_860_43_n_16,
     sub_860_43_n_17, sub_860_43_n_18, sub_860_43_n_19, sub_860_43_n_20,
     sub_860_43_n_21, sub_860_43_n_22, sub_860_43_n_23, sub_860_43_n_24,
     sub_860_43_n_25, sub_860_43_n_26, sub_860_43_n_27, sub_860_43_n_28,
     sub_860_43_n_29, sub_860_43_n_30, sub_860_43_n_31, sub_860_43_n_32,
     sub_860_43_n_33, sub_860_43_n_34, sub_860_43_n_35, sub_860_43_n_37,
     sub_860_43_n_38, sub_860_43_n_39, sub_860_43_n_40, sub_860_43_n_41,
     sub_860_43_n_42, sub_860_43_n_43, sub_860_43_n_44, sub_860_43_n_46,
     sub_860_43_n_47, sub_860_43_n_48, sub_860_43_n_49, sub_860_43_n_50,
     sub_860_43_n_51, sub_860_43_n_52, sub_860_43_n_53, sub_860_43_n_54,
     sub_860_43_n_55, sub_860_43_n_56, sub_860_43_n_57, sub_860_43_n_58,
     sub_860_43_n_59, sub_860_43_n_60, sub_860_43_n_61, sub_860_43_n_62,
     sub_860_43_n_63, sub_860_43_n_64, sub_860_43_n_65, sub_860_43_n_66,
     sub_860_43_n_67, sub_860_43_n_68, sub_860_43_n_69, sub_860_43_n_70,
     sub_860_43_n_71, sub_860_43_n_72, sub_860_43_n_73, sub_860_43_n_74,
     sub_860_43_n_75, sub_860_43_n_76, sub_860_43_n_77, sub_860_43_n_78,
     sub_860_43_n_79, sub_860_43_n_80, sub_860_43_n_81, sub_860_43_n_82,
     sub_860_43_n_83, sub_860_43_n_84, sub_860_43_n_85, sub_860_43_n_87,
     sub_860_43_n_88, sub_860_43_n_89, sub_860_43_n_90, sub_860_43_n_91,
     sub_860_43_n_92, sub_860_43_n_93, sub_860_43_n_94, sub_860_43_n_95,
     sub_860_43_n_96, sub_860_43_n_97, sub_860_43_n_98, sub_860_43_n_99,
     sub_860_43_n_100, sub_860_43_n_101, sub_860_43_n_102, sub_860_43_n_103,
     sub_860_43_n_104, sub_860_43_n_105, sub_860_43_n_106, sub_860_43_n_107,
     sub_860_43_n_108, sub_860_43_n_109, sub_860_43_n_110, sub_860_43_n_111,
     sub_860_43_n_112, sub_860_43_n_113, sub_860_43_n_114, sub_860_43_n_115,
     sub_860_43_n_116, sub_860_43_n_117, sub_860_43_n_118, sub_860_43_n_119,
     sub_860_43_n_120, sub_860_43_n_121, sub_860_43_n_122, sub_860_43_n_123,
     sub_860_43_n_124, sub_860_43_n_125, sub_860_43_n_126, sub_860_43_n_127,
     sub_860_43_n_128, sub_860_43_n_129, sub_860_43_n_130, sub_860_43_n_131,
     sub_860_43_n_133, sub_860_43_n_134, sub_860_43_n_135, sub_860_43_n_136,
     sub_860_43_n_137, sub_860_43_n_139, sub_860_43_n_140, sub_860_43_n_141,
     sub_860_43_n_142, sub_860_43_n_145, sub_860_43_n_146, sub_860_43_n_147,
     sub_860_43_n_148, sub_860_43_n_149, sub_860_43_n_150, sub_860_43_n_154,
     sub_860_43_n_155, sub_860_43_n_156, sub_860_43_n_157, sub_860_43_n_158,
     sub_860_43_n_163, sub_860_43_n_165, sub_860_43_n_166, sub_860_43_n_167,
     sub_860_43_n_168, sub_860_43_n_169, sub_860_43_n_176, sub_890_40_n_0,
     sub_890_40_n_1, sub_890_40_n_2, sub_890_40_n_3, sub_890_40_n_4,
     sub_890_40_n_5, sub_890_40_n_6, sub_890_40_n_7, sub_890_40_n_8,
     sub_890_40_n_9, sub_890_40_n_10, sub_890_40_n_11, sub_890_40_n_12,
     sub_890_40_n_13, sub_890_40_n_14, sub_890_40_n_15, sub_890_40_n_16,
     sub_890_40_n_17, sub_890_40_n_18, sub_890_40_n_19, sub_890_40_n_20,
     sub_890_40_n_21, sub_890_40_n_22, sub_890_40_n_23, sub_890_40_n_24,
     sub_890_40_n_25, sub_890_40_n_26, sub_890_40_n_27, sub_890_40_n_28,
     sub_890_40_n_30, sub_890_40_n_31, sub_890_40_n_32, sub_890_40_n_33,
     sub_890_40_n_34, sub_890_40_n_35, sub_890_40_n_36, sub_890_40_n_37,
     sub_890_40_n_38, sub_890_40_n_40, sub_890_40_n_41, sub_890_40_n_42,
     sub_890_40_n_43, sub_890_40_n_45, sub_890_40_n_46, sub_890_40_n_47,
     sub_890_40_n_48, sub_890_40_n_49, sub_890_40_n_50, sub_890_40_n_51,
     sub_890_40_n_52, sub_890_40_n_53, sub_890_40_n_54, sub_890_40_n_55,
     sub_890_40_n_56, sub_890_40_n_57, sub_890_40_n_58, sub_890_40_n_59,
     sub_890_40_n_60, sub_890_40_n_61, sub_890_40_n_62, sub_890_40_n_63,
     sub_890_40_n_64, sub_890_40_n_65, sub_890_40_n_66, sub_890_40_n_67,
     sub_890_40_n_68, sub_890_40_n_69, sub_890_40_n_70, sub_890_40_n_71,
     sub_890_40_n_72, sub_890_40_n_73, sub_890_40_n_74, sub_890_40_n_75,
     sub_890_40_n_76, sub_890_40_n_77, sub_890_40_n_78, sub_890_40_n_79,
     sub_890_40_n_80, sub_890_40_n_81, sub_890_40_n_82, sub_890_40_n_83,
     sub_890_40_n_84, sub_890_40_n_85, sub_890_40_n_86, sub_890_40_n_87,
     sub_890_40_n_88, sub_890_40_n_89, sub_890_40_n_90, sub_890_40_n_91,
     sub_890_40_n_92, sub_890_40_n_94, sub_890_40_n_95, sub_890_40_n_96,
     sub_890_40_n_97, sub_890_40_n_98, sub_890_40_n_99, sub_890_40_n_100,
     sub_890_40_n_101, sub_890_40_n_102, sub_890_40_n_103, sub_890_40_n_104,
     sub_890_40_n_105, sub_890_40_n_106, sub_890_40_n_107, sub_890_40_n_108,
     sub_890_40_n_109, sub_890_40_n_110, sub_890_40_n_111, sub_890_40_n_112,
     sub_890_40_n_113, sub_890_40_n_114, sub_890_40_n_115, sub_890_40_n_116,
     sub_890_40_n_117, sub_890_40_n_118, sub_890_40_n_119, sub_890_40_n_120,
     sub_890_40_n_121, sub_890_40_n_122, sub_890_40_n_123, sub_890_40_n_124,
     sub_890_40_n_125, sub_890_40_n_126, sub_890_40_n_127, sub_890_40_n_128,
     sub_890_40_n_129, sub_890_40_n_130, sub_890_40_n_131, sub_890_40_n_132,
     sub_890_40_n_133, sub_890_40_n_134, sub_890_40_n_135, sub_890_40_n_136,
     sub_890_40_n_137, sub_890_40_n_138, sub_890_40_n_139, sub_890_40_n_140,
     sub_890_40_n_141, sub_890_40_n_142, sub_890_40_n_143, sub_890_40_n_144,
     sub_890_40_n_145, sub_890_40_n_146, sub_890_40_n_147, sub_890_40_n_149,
     sub_890_40_n_150, sub_890_40_n_151, sub_890_40_n_152, sub_890_40_n_153,
     sub_890_40_n_155, sub_890_40_n_156, sub_890_40_n_157, sub_890_40_n_158,
     sub_890_40_n_161, sub_890_40_n_162, sub_890_40_n_163, sub_890_40_n_164,
     sub_890_40_n_167, sub_890_40_n_168, sub_890_40_n_169, sub_890_40_n_170,
     sub_890_40_n_171, sub_890_40_n_172, sub_890_40_n_173, sub_890_40_n_179,
     sub_890_40_n_180, sub_890_40_n_181, sub_890_40_n_182, sub_890_40_n_183,
     sub_890_40_n_184, sub_890_40_n_191, sub_890_40_n_192, sub_920_38_n_0,
     sub_920_38_n_1, sub_920_38_n_2, sub_920_38_n_3, sub_920_38_n_4,
     sub_920_38_n_5, sub_920_38_n_6, sub_920_38_n_7, sub_920_38_n_8,
     sub_920_38_n_9, sub_920_38_n_10, sub_920_38_n_11, sub_920_38_n_12,
     sub_920_38_n_13, sub_920_38_n_14, sub_920_38_n_15, sub_920_38_n_16,
     sub_920_38_n_17, sub_920_38_n_18, sub_920_38_n_19, sub_920_38_n_20,
     sub_920_38_n_21, sub_920_38_n_22, sub_920_38_n_23, sub_920_38_n_24,
     sub_920_38_n_25, sub_920_38_n_26, sub_920_38_n_27, sub_920_38_n_28,
     sub_920_38_n_29, sub_920_38_n_30, sub_920_38_n_31, sub_920_38_n_32,
     sub_920_38_n_33, sub_920_38_n_34, sub_920_38_n_35, sub_920_38_n_36,
     sub_920_38_n_37, sub_920_38_n_38, sub_920_38_n_39, sub_920_38_n_40,
     sub_920_38_n_41, sub_920_38_n_42, sub_920_38_n_44, sub_920_38_n_45,
     sub_920_38_n_46, sub_920_38_n_47, sub_920_38_n_48, sub_920_38_n_49,
     sub_920_38_n_50, sub_920_38_n_51, sub_920_38_n_52, sub_920_38_n_53,
     sub_920_38_n_54, sub_920_38_n_55, sub_920_38_n_56, sub_920_38_n_57,
     sub_920_38_n_58, sub_920_38_n_59, sub_920_38_n_60, sub_920_38_n_61,
     sub_920_38_n_62, sub_920_38_n_63, sub_920_38_n_64, sub_920_38_n_65,
     sub_920_38_n_66, sub_920_38_n_67, sub_920_38_n_68, sub_920_38_n_69,
     sub_920_38_n_70, sub_920_38_n_71, sub_920_38_n_72, sub_920_38_n_73,
     sub_920_38_n_74, sub_920_38_n_75, sub_920_38_n_76, sub_920_38_n_77,
     sub_920_38_n_78, sub_920_38_n_79, sub_920_38_n_80, sub_920_38_n_81,
     sub_920_38_n_82, sub_920_38_n_83, sub_920_38_n_84, sub_920_38_n_85,
     sub_920_38_n_86, sub_920_38_n_87, sub_920_38_n_88, sub_920_38_n_89,
     sub_920_38_n_90, sub_920_38_n_91, sub_920_38_n_92, sub_920_38_n_93,
     sub_920_38_n_94, sub_920_38_n_95, sub_920_38_n_96, sub_920_38_n_97,
     sub_920_38_n_98, sub_920_38_n_99, sub_920_38_n_100, sub_920_38_n_102,
     sub_920_38_n_103, sub_920_38_n_104, sub_920_38_n_105, sub_920_38_n_106,
     sub_920_38_n_107, sub_920_38_n_108, sub_920_38_n_109, sub_920_38_n_110,
     sub_920_38_n_111, sub_920_38_n_112, sub_920_38_n_113, sub_920_38_n_114,
     sub_920_38_n_115, sub_920_38_n_116, sub_920_38_n_117, sub_920_38_n_118,
     sub_920_38_n_119, sub_920_38_n_120, sub_920_38_n_121, sub_920_38_n_122,
     sub_920_38_n_123, sub_920_38_n_124, sub_920_38_n_125, sub_920_38_n_126,
     sub_920_38_n_127, sub_920_38_n_128, sub_920_38_n_129, sub_920_38_n_130,
     sub_920_38_n_131, sub_920_38_n_132, sub_920_38_n_133, sub_920_38_n_134,
     sub_920_38_n_135, sub_920_38_n_136, sub_920_38_n_137, sub_920_38_n_138,
     sub_920_38_n_139, sub_920_38_n_140, sub_920_38_n_141, sub_920_38_n_142,
     sub_920_38_n_143, sub_920_38_n_144, sub_920_38_n_145, sub_920_38_n_146,
     sub_920_38_n_147, sub_920_38_n_148, sub_920_38_n_149, sub_920_38_n_150,
     sub_920_38_n_151, sub_920_38_n_152, sub_920_38_n_153, sub_920_38_n_154,
     sub_920_38_n_155, sub_920_38_n_156, sub_920_38_n_157, sub_920_38_n_158,
     sub_920_38_n_159, sub_920_38_n_161, sub_920_38_n_162, sub_920_38_n_163,
     sub_920_38_n_164, sub_920_38_n_165, sub_920_38_n_166, sub_920_38_n_167,
     sub_920_38_n_168, sub_920_38_n_170, sub_920_38_n_171, sub_920_38_n_172,
     sub_920_38_n_173, sub_920_38_n_176, sub_920_38_n_177, sub_920_38_n_178,
     sub_920_38_n_179, sub_920_38_n_180, sub_920_38_n_184, sub_920_38_n_185,
     sub_920_38_n_186, sub_920_38_n_187, sub_920_38_n_188, sub_920_38_n_189,
     sub_920_38_n_190, sub_920_38_n_196, sub_920_38_n_197, sub_920_38_n_198,
     sub_920_38_n_199, sub_920_38_n_200, sub_920_38_n_201, sub_920_38_n_202,
     sub_920_38_n_203, sub_920_38_n_204, sub_920_38_n_212, sub_920_38_n_213,
     sub_920_38_n_215, sub_950_37_n_0, sub_950_37_n_1, sub_950_37_n_2,
     sub_950_37_n_3, sub_950_37_n_4, sub_950_37_n_5, sub_950_37_n_6,
     sub_950_37_n_7, sub_950_37_n_8, sub_950_37_n_9, sub_950_37_n_10,
     sub_950_37_n_11, sub_950_37_n_12, sub_950_37_n_13, sub_950_37_n_14,
     sub_950_37_n_15, sub_950_37_n_16, sub_950_37_n_17, sub_950_37_n_18,
     sub_950_37_n_19, sub_950_37_n_20, sub_950_37_n_21, sub_950_37_n_22,
     sub_950_37_n_23, sub_950_37_n_24, sub_950_37_n_25, sub_950_37_n_26,
     sub_950_37_n_27, sub_950_37_n_28, sub_950_37_n_29, sub_950_37_n_30,
     sub_950_37_n_31, sub_950_37_n_32, sub_950_37_n_33, sub_950_37_n_34,
     sub_950_37_n_35, sub_950_37_n_36, sub_950_37_n_37, sub_950_37_n_38,
     sub_950_37_n_39, sub_950_37_n_40, sub_950_37_n_41, sub_950_37_n_42,
     sub_950_37_n_43, sub_950_37_n_44, sub_950_37_n_45, sub_950_37_n_46,
     sub_950_37_n_47, sub_950_37_n_48, sub_950_37_n_49, sub_950_37_n_51,
     sub_950_37_n_52, sub_950_37_n_53, sub_950_37_n_54, sub_950_37_n_55,
     sub_950_37_n_56, sub_950_37_n_57, sub_950_37_n_58, sub_950_37_n_59,
     sub_950_37_n_61, sub_950_37_n_62, sub_950_37_n_63, sub_950_37_n_64,
     sub_950_37_n_65, sub_950_37_n_66, sub_950_37_n_67, sub_950_37_n_68,
     sub_950_37_n_69, sub_950_37_n_70, sub_950_37_n_71, sub_950_37_n_72,
     sub_950_37_n_73, sub_950_37_n_74, sub_950_37_n_75, sub_950_37_n_76,
     sub_950_37_n_77, sub_950_37_n_78, sub_950_37_n_79, sub_950_37_n_80,
     sub_950_37_n_81, sub_950_37_n_82, sub_950_37_n_83, sub_950_37_n_84,
     sub_950_37_n_85, sub_950_37_n_86, sub_950_37_n_87, sub_950_37_n_88,
     sub_950_37_n_89, sub_950_37_n_90, sub_950_37_n_91, sub_950_37_n_92,
     sub_950_37_n_93, sub_950_37_n_94, sub_950_37_n_95, sub_950_37_n_96,
     sub_950_37_n_97, sub_950_37_n_98, sub_950_37_n_100, sub_950_37_n_101,
     sub_950_37_n_102, sub_950_37_n_103, sub_950_37_n_104, sub_950_37_n_105,
     sub_950_37_n_106, sub_950_37_n_107, sub_950_37_n_108, sub_950_37_n_109,
     sub_950_37_n_110, sub_950_37_n_111, sub_950_37_n_112, sub_950_37_n_113,
     sub_950_37_n_114, sub_950_37_n_115, sub_950_37_n_116, sub_950_37_n_117,
     sub_950_37_n_118, sub_950_37_n_119, sub_950_37_n_120, sub_950_37_n_121,
     sub_950_37_n_122, sub_950_37_n_123, sub_950_37_n_124, sub_950_37_n_125,
     sub_950_37_n_126, sub_950_37_n_127, sub_950_37_n_128, sub_950_37_n_129,
     sub_950_37_n_130, sub_950_37_n_131, sub_950_37_n_132, sub_950_37_n_133,
     sub_950_37_n_134, sub_950_37_n_135, sub_950_37_n_136, sub_950_37_n_137,
     sub_950_37_n_138, sub_950_37_n_139, sub_950_37_n_140, sub_950_37_n_141,
     sub_950_37_n_142, sub_950_37_n_143, sub_950_37_n_144, sub_950_37_n_145,
     sub_950_37_n_146, sub_950_37_n_147, sub_950_37_n_149, sub_950_37_n_150,
     sub_950_37_n_151, sub_950_37_n_152, sub_950_37_n_153, sub_950_37_n_155,
     sub_950_37_n_156, sub_950_37_n_157, sub_950_37_n_158, sub_950_37_n_159,
     sub_950_37_n_161, sub_950_37_n_162, sub_950_37_n_163, sub_950_37_n_164,
     sub_950_37_n_165, sub_950_37_n_169, sub_950_37_n_170, sub_950_37_n_171,
     sub_950_37_n_172, sub_950_37_n_173, sub_950_37_n_174, sub_950_37_n_175,
     sub_950_37_n_176, sub_950_37_n_177, sub_950_37_n_178, sub_950_37_n_184,
     sub_950_37_n_185, sub_950_37_n_187, sub_950_37_n_188, sub_950_37_n_189,
     sub_950_37_n_190, sub_950_37_n_191, sub_950_37_n_192, sub_950_37_n_193,
     sub_950_37_n_201, sub_950_37_n_202, sub_950_37_n_203, sub_980_36_n_0,
     sub_980_36_n_1, sub_980_36_n_2, sub_980_36_n_3, sub_980_36_n_4,
     sub_980_36_n_5, sub_980_36_n_6, sub_980_36_n_7, sub_980_36_n_8,
     sub_980_36_n_9, sub_980_36_n_10, sub_980_36_n_11, sub_980_36_n_12,
     sub_980_36_n_13, sub_980_36_n_14, sub_980_36_n_15, sub_980_36_n_16,
     sub_980_36_n_17, sub_980_36_n_18, sub_980_36_n_19, sub_980_36_n_20,
     sub_980_36_n_21, sub_980_36_n_22, sub_980_36_n_23, sub_980_36_n_24,
     sub_980_36_n_25, sub_980_36_n_26, sub_980_36_n_27, sub_980_36_n_28,
     sub_980_36_n_29, sub_980_36_n_30, sub_980_36_n_31, sub_980_36_n_32,
     sub_980_36_n_33, sub_980_36_n_34, sub_980_36_n_35, sub_980_36_n_36,
     sub_980_36_n_37, sub_980_36_n_38, sub_980_36_n_39, sub_980_36_n_40,
     sub_980_36_n_41, sub_980_36_n_42, sub_980_36_n_43, sub_980_36_n_44,
     sub_980_36_n_45, sub_980_36_n_46, sub_980_36_n_47, sub_980_36_n_48,
     sub_980_36_n_50, sub_980_36_n_51, sub_980_36_n_52, sub_980_36_n_53,
     sub_980_36_n_54, sub_980_36_n_55, sub_980_36_n_56, sub_980_36_n_57,
     sub_980_36_n_58, sub_980_36_n_59, sub_980_36_n_60, sub_980_36_n_61,
     sub_980_36_n_62, sub_980_36_n_63, sub_980_36_n_64, sub_980_36_n_65,
     sub_980_36_n_66, sub_980_36_n_67, sub_980_36_n_68, sub_980_36_n_69,
     sub_980_36_n_70, sub_980_36_n_71, sub_980_36_n_72, sub_980_36_n_73,
     sub_980_36_n_74, sub_980_36_n_75, sub_980_36_n_76, sub_980_36_n_77,
     sub_980_36_n_78, sub_980_36_n_79, sub_980_36_n_80, sub_980_36_n_81,
     sub_980_36_n_82, sub_980_36_n_83, sub_980_36_n_84, sub_980_36_n_85,
     sub_980_36_n_86, sub_980_36_n_87, sub_980_36_n_88, sub_980_36_n_89,
     sub_980_36_n_90, sub_980_36_n_91, sub_980_36_n_92, sub_980_36_n_93,
     sub_980_36_n_94, sub_980_36_n_95, sub_980_36_n_96, sub_980_36_n_97,
     sub_980_36_n_98, sub_980_36_n_99, sub_980_36_n_100, sub_980_36_n_101,
     sub_980_36_n_102, sub_980_36_n_103, sub_980_36_n_104, sub_980_36_n_105,
     sub_980_36_n_106, sub_980_36_n_107, sub_980_36_n_108, sub_980_36_n_109,
     sub_980_36_n_110, sub_980_36_n_111, sub_980_36_n_112, sub_980_36_n_113,
     sub_980_36_n_114, sub_980_36_n_115, sub_980_36_n_116, sub_980_36_n_118,
     sub_980_36_n_119, sub_980_36_n_120, sub_980_36_n_121, sub_980_36_n_122,
     sub_980_36_n_123, sub_980_36_n_124, sub_980_36_n_125, sub_980_36_n_126,
     sub_980_36_n_127, sub_980_36_n_128, sub_980_36_n_129, sub_980_36_n_130,
     sub_980_36_n_131, sub_980_36_n_132, sub_980_36_n_133, sub_980_36_n_134,
     sub_980_36_n_135, sub_980_36_n_136, sub_980_36_n_137, sub_980_36_n_138,
     sub_980_36_n_139, sub_980_36_n_140, sub_980_36_n_141, sub_980_36_n_142,
     sub_980_36_n_143, sub_980_36_n_144, sub_980_36_n_145, sub_980_36_n_146,
     sub_980_36_n_147, sub_980_36_n_148, sub_980_36_n_149, sub_980_36_n_150,
     sub_980_36_n_151, sub_980_36_n_152, sub_980_36_n_153, sub_980_36_n_154,
     sub_980_36_n_155, sub_980_36_n_156, sub_980_36_n_157, sub_980_36_n_158,
     sub_980_36_n_159, sub_980_36_n_160, sub_980_36_n_161, sub_980_36_n_162,
     sub_980_36_n_163, sub_980_36_n_164, sub_980_36_n_166, sub_980_36_n_167,
     sub_980_36_n_168, sub_980_36_n_169, sub_980_36_n_170, sub_980_36_n_171,
     sub_980_36_n_172, sub_980_36_n_173, sub_980_36_n_174, sub_980_36_n_175,
     sub_980_36_n_176, sub_980_36_n_177, sub_980_36_n_179, sub_980_36_n_180,
     sub_980_36_n_181, sub_980_36_n_182, sub_980_36_n_185, sub_980_36_n_186,
     sub_980_36_n_187, sub_980_36_n_188, sub_980_36_n_189, sub_980_36_n_193,
     sub_980_36_n_194, sub_980_36_n_195, sub_980_36_n_196, sub_980_36_n_197,
     sub_980_36_n_198, sub_980_36_n_199, sub_980_36_n_200, sub_980_36_n_201,
     sub_980_36_n_207, sub_980_36_n_208, sub_980_36_n_209, sub_980_36_n_211,
     sub_980_36_n_212, sub_980_36_n_213, sub_980_36_n_214, sub_980_36_n_215,
     sub_980_36_n_224, sub_980_36_n_225, sub_980_36_n_226, sub_980_36_n_227,
     sub_1010_35_n_0, sub_1010_35_n_1, sub_1010_35_n_2, sub_1010_35_n_3,
     sub_1010_35_n_4, sub_1010_35_n_5, sub_1010_35_n_6, sub_1010_35_n_7,
     sub_1010_35_n_8, sub_1010_35_n_9, sub_1010_35_n_10, sub_1010_35_n_11,
     sub_1010_35_n_12, sub_1010_35_n_13, sub_1010_35_n_14, sub_1010_35_n_15,
     sub_1010_35_n_16, sub_1010_35_n_17, sub_1010_35_n_18, sub_1010_35_n_19,
     sub_1010_35_n_20, sub_1010_35_n_21, sub_1010_35_n_22, sub_1010_35_n_23,
     sub_1010_35_n_24, sub_1010_35_n_25, sub_1010_35_n_26, sub_1010_35_n_27,
     sub_1010_35_n_28, sub_1010_35_n_29, sub_1010_35_n_30, sub_1010_35_n_31,
     sub_1010_35_n_32, sub_1010_35_n_33, sub_1010_35_n_34, sub_1010_35_n_35,
     sub_1010_35_n_36, sub_1010_35_n_37, sub_1010_35_n_38, sub_1010_35_n_39,
     sub_1010_35_n_40, sub_1010_35_n_41, sub_1010_35_n_42, sub_1010_35_n_43,
     sub_1010_35_n_44, sub_1010_35_n_45, sub_1010_35_n_46, sub_1010_35_n_47,
     sub_1010_35_n_49, sub_1010_35_n_50, sub_1010_35_n_51, sub_1010_35_n_52,
     sub_1010_35_n_53, sub_1010_35_n_54, sub_1010_35_n_55, sub_1010_35_n_56,
     sub_1010_35_n_57, sub_1010_35_n_58, sub_1010_35_n_59, sub_1010_35_n_60,
     sub_1010_35_n_61, sub_1010_35_n_62, sub_1010_35_n_63, sub_1010_35_n_64,
     sub_1010_35_n_65, sub_1010_35_n_66, sub_1010_35_n_67, sub_1010_35_n_68,
     sub_1010_35_n_69, sub_1010_35_n_70, sub_1010_35_n_71, sub_1010_35_n_72,
     sub_1010_35_n_73, sub_1010_35_n_74, sub_1010_35_n_75, sub_1010_35_n_76,
     sub_1010_35_n_77, sub_1010_35_n_78, sub_1010_35_n_79, sub_1010_35_n_80,
     sub_1010_35_n_81, sub_1010_35_n_82, sub_1010_35_n_83, sub_1010_35_n_84,
     sub_1010_35_n_85, sub_1010_35_n_86, sub_1010_35_n_87, sub_1010_35_n_88,
     sub_1010_35_n_89, sub_1010_35_n_90, sub_1010_35_n_91, sub_1010_35_n_92,
     sub_1010_35_n_93, sub_1010_35_n_94, sub_1010_35_n_95, sub_1010_35_n_96,
     sub_1010_35_n_97, sub_1010_35_n_98, sub_1010_35_n_99, sub_1010_35_n_100,
     sub_1010_35_n_101, sub_1010_35_n_103, sub_1010_35_n_104, sub_1010_35_n_105,
     sub_1010_35_n_106, sub_1010_35_n_107, sub_1010_35_n_108, sub_1010_35_n_109,
     sub_1010_35_n_110, sub_1010_35_n_111, sub_1010_35_n_112, sub_1010_35_n_113,
     sub_1010_35_n_114, sub_1010_35_n_115, sub_1010_35_n_116, sub_1010_35_n_117,
     sub_1010_35_n_118, sub_1010_35_n_119, sub_1010_35_n_120, sub_1010_35_n_121,
     sub_1010_35_n_122, sub_1010_35_n_123, sub_1010_35_n_124, sub_1010_35_n_125,
     sub_1010_35_n_126, sub_1010_35_n_127, sub_1010_35_n_128, sub_1010_35_n_129,
     sub_1010_35_n_130, sub_1010_35_n_131, sub_1010_35_n_132, sub_1010_35_n_133,
     sub_1010_35_n_134, sub_1010_35_n_135, sub_1010_35_n_136, sub_1010_35_n_137,
     sub_1010_35_n_138, sub_1010_35_n_139, sub_1010_35_n_140, sub_1010_35_n_141,
     sub_1010_35_n_142, sub_1010_35_n_143, sub_1010_35_n_144, sub_1010_35_n_145,
     sub_1010_35_n_146, sub_1010_35_n_147, sub_1010_35_n_148, sub_1010_35_n_149,
     sub_1010_35_n_150, sub_1010_35_n_151, sub_1010_35_n_152, sub_1010_35_n_153,
     sub_1010_35_n_154, sub_1010_35_n_155, sub_1010_35_n_156, sub_1010_35_n_157,
     sub_1010_35_n_158, sub_1010_35_n_159, sub_1010_35_n_160, sub_1010_35_n_161,
     sub_1010_35_n_162, sub_1010_35_n_163, sub_1010_35_n_164, sub_1010_35_n_165,
     sub_1010_35_n_166, sub_1010_35_n_167, sub_1010_35_n_168, sub_1010_35_n_169,
     sub_1010_35_n_170, sub_1010_35_n_171, sub_1010_35_n_172, sub_1010_35_n_174,
     sub_1010_35_n_175, sub_1010_35_n_176, sub_1010_35_n_177, sub_1010_35_n_178,
     sub_1010_35_n_179, sub_1010_35_n_180, sub_1010_35_n_181, sub_1010_35_n_182,
     sub_1010_35_n_183, sub_1010_35_n_184, sub_1010_35_n_186, sub_1010_35_n_187,
     sub_1010_35_n_188, sub_1010_35_n_189, sub_1010_35_n_192, sub_1010_35_n_193,
     sub_1010_35_n_194, sub_1010_35_n_195, sub_1010_35_n_196, sub_1010_35_n_197,
     sub_1010_35_n_201, sub_1010_35_n_202, sub_1010_35_n_203, sub_1010_35_n_204,
     sub_1010_35_n_205, sub_1010_35_n_206, sub_1010_35_n_207, sub_1010_35_n_208,
     sub_1010_35_n_209, sub_1010_35_n_210, sub_1010_35_n_211, sub_1010_35_n_217,
     sub_1010_35_n_219, sub_1010_35_n_220, sub_1010_35_n_221, sub_1010_35_n_222,
     sub_1010_35_n_231, sub_1010_35_n_232, sub_1010_35_n_233, sub_1010_35_n_234,
     sub_1040_34_n_0, sub_1040_34_n_1, sub_1040_34_n_2, sub_1040_34_n_3,
     sub_1040_34_n_4, sub_1040_34_n_5, sub_1040_34_n_6, sub_1040_34_n_7,
     sub_1040_34_n_8, sub_1040_34_n_9, sub_1040_34_n_10, sub_1040_34_n_11,
     sub_1040_34_n_12, sub_1040_34_n_13, sub_1040_34_n_14, sub_1040_34_n_15,
     sub_1040_34_n_16, sub_1040_34_n_17, sub_1040_34_n_18, sub_1040_34_n_19,
     sub_1040_34_n_20, sub_1040_34_n_21, sub_1040_34_n_22, sub_1040_34_n_23,
     sub_1040_34_n_24, sub_1040_34_n_25, sub_1040_34_n_26, sub_1040_34_n_27,
     sub_1040_34_n_28, sub_1040_34_n_29, sub_1040_34_n_30, sub_1040_34_n_31,
     sub_1040_34_n_32, sub_1040_34_n_33, sub_1040_34_n_34, sub_1040_34_n_35,
     sub_1040_34_n_36, sub_1040_34_n_37, sub_1040_34_n_38, sub_1040_34_n_39,
     sub_1040_34_n_40, sub_1040_34_n_41, sub_1040_34_n_42, sub_1040_34_n_44,
     sub_1040_34_n_45, sub_1040_34_n_46, sub_1040_34_n_47, sub_1040_34_n_48,
     sub_1040_34_n_49, sub_1040_34_n_50, sub_1040_34_n_52, sub_1040_34_n_53,
     sub_1040_34_n_54, sub_1040_34_n_55, sub_1040_34_n_56, sub_1040_34_n_57,
     sub_1040_34_n_58, sub_1040_34_n_59, sub_1040_34_n_60, sub_1040_34_n_61,
     sub_1040_34_n_62, sub_1040_34_n_63, sub_1040_34_n_64, sub_1040_34_n_65,
     sub_1040_34_n_66, sub_1040_34_n_67, sub_1040_34_n_68, sub_1040_34_n_69,
     sub_1040_34_n_70, sub_1040_34_n_71, sub_1040_34_n_72, sub_1040_34_n_73,
     sub_1040_34_n_74, sub_1040_34_n_75, sub_1040_34_n_76, sub_1040_34_n_77,
     sub_1040_34_n_78, sub_1040_34_n_79, sub_1040_34_n_80, sub_1040_34_n_81,
     sub_1040_34_n_82, sub_1040_34_n_83, sub_1040_34_n_84, sub_1040_34_n_85,
     sub_1040_34_n_86, sub_1040_34_n_87, sub_1040_34_n_88, sub_1040_34_n_89,
     sub_1040_34_n_90, sub_1040_34_n_91, sub_1040_34_n_92, sub_1040_34_n_93,
     sub_1040_34_n_94, sub_1040_34_n_95, sub_1040_34_n_96, sub_1040_34_n_97,
     sub_1040_34_n_98, sub_1040_34_n_99, sub_1040_34_n_100, sub_1040_34_n_101,
     sub_1040_34_n_102, sub_1040_34_n_103, sub_1040_34_n_104, sub_1040_34_n_105,
     sub_1040_34_n_106, sub_1040_34_n_107, sub_1040_34_n_108, sub_1040_34_n_109,
     sub_1040_34_n_110, sub_1040_34_n_111, sub_1040_34_n_113, sub_1040_34_n_114,
     sub_1040_34_n_115, sub_1040_34_n_116, sub_1040_34_n_117, sub_1040_34_n_118,
     sub_1040_34_n_119, sub_1040_34_n_120, sub_1040_34_n_121, sub_1040_34_n_122,
     sub_1040_34_n_123, sub_1040_34_n_124, sub_1040_34_n_125, sub_1040_34_n_126,
     sub_1040_34_n_127, sub_1040_34_n_128, sub_1040_34_n_129, sub_1040_34_n_130,
     sub_1040_34_n_131, sub_1040_34_n_132, sub_1040_34_n_133, sub_1040_34_n_134,
     sub_1040_34_n_135, sub_1040_34_n_136, sub_1040_34_n_137, sub_1040_34_n_138,
     sub_1040_34_n_139, sub_1040_34_n_140, sub_1040_34_n_141, sub_1040_34_n_142,
     sub_1040_34_n_143, sub_1040_34_n_144, sub_1040_34_n_145, sub_1040_34_n_146,
     sub_1040_34_n_147, sub_1040_34_n_148, sub_1040_34_n_149, sub_1040_34_n_150,
     sub_1040_34_n_151, sub_1040_34_n_152, sub_1040_34_n_153, sub_1040_34_n_154,
     sub_1040_34_n_155, sub_1040_34_n_156, sub_1040_34_n_157, sub_1040_34_n_158,
     sub_1040_34_n_159, sub_1040_34_n_160, sub_1040_34_n_161, sub_1040_34_n_162,
     sub_1040_34_n_163, sub_1040_34_n_164, sub_1040_34_n_165, sub_1040_34_n_166,
     sub_1040_34_n_167, sub_1040_34_n_168, sub_1040_34_n_169, sub_1040_34_n_170,
     sub_1040_34_n_171, sub_1040_34_n_173, sub_1040_34_n_174, sub_1040_34_n_175,
     sub_1040_34_n_176, sub_1040_34_n_177, sub_1040_34_n_178, sub_1040_34_n_179,
     sub_1040_34_n_180, sub_1040_34_n_182, sub_1040_34_n_183, sub_1040_34_n_184,
     sub_1040_34_n_185, sub_1040_34_n_188, sub_1040_34_n_189, sub_1040_34_n_190,
     sub_1040_34_n_191, sub_1040_34_n_192, sub_1040_34_n_193, sub_1040_34_n_194,
     sub_1040_34_n_197, sub_1040_34_n_198, sub_1040_34_n_199, sub_1040_34_n_200,
     sub_1040_34_n_201, sub_1040_34_n_202, sub_1040_34_n_203, sub_1040_34_n_204,
     sub_1040_34_n_205, sub_1040_34_n_206, sub_1040_34_n_212, sub_1040_34_n_214,
     sub_1040_34_n_215, sub_1040_34_n_216, sub_1040_34_n_217, sub_1040_34_n_218,
     sub_1040_34_n_219, sub_1040_34_n_228, sub_1040_34_n_229, sub_1040_34_n_230,
     sub_1040_34_n_231, sub_1040_34_n_232, sub_1070_33_n_0, sub_1070_33_n_1,
     sub_1070_33_n_2, sub_1070_33_n_3, sub_1070_33_n_4, sub_1070_33_n_5,
     sub_1070_33_n_6, sub_1070_33_n_7, sub_1070_33_n_8, sub_1070_33_n_9,
     sub_1070_33_n_10, sub_1070_33_n_11, sub_1070_33_n_12, sub_1070_33_n_13,
     sub_1070_33_n_14, sub_1070_33_n_15, sub_1070_33_n_16, sub_1070_33_n_17,
     sub_1070_33_n_18, sub_1070_33_n_19, sub_1070_33_n_20, sub_1070_33_n_21,
     sub_1070_33_n_22, sub_1070_33_n_23, sub_1070_33_n_24, sub_1070_33_n_25,
     sub_1070_33_n_26, sub_1070_33_n_27, sub_1070_33_n_28, sub_1070_33_n_29,
     sub_1070_33_n_30, sub_1070_33_n_31, sub_1070_33_n_32, sub_1070_33_n_33,
     sub_1070_33_n_34, sub_1070_33_n_35, sub_1070_33_n_36, sub_1070_33_n_37,
     sub_1070_33_n_38, sub_1070_33_n_39, sub_1070_33_n_40, sub_1070_33_n_41,
     sub_1070_33_n_42, sub_1070_33_n_43, sub_1070_33_n_45, sub_1070_33_n_46,
     sub_1070_33_n_47, sub_1070_33_n_48, sub_1070_33_n_49, sub_1070_33_n_50,
     sub_1070_33_n_51, sub_1070_33_n_52, sub_1070_33_n_53, sub_1070_33_n_54,
     sub_1070_33_n_56, sub_1070_33_n_57, sub_1070_33_n_58, sub_1070_33_n_59,
     sub_1070_33_n_60, sub_1070_33_n_61, sub_1070_33_n_62, sub_1070_33_n_63,
     sub_1070_33_n_64, sub_1070_33_n_65, sub_1070_33_n_66, sub_1070_33_n_67,
     sub_1070_33_n_68, sub_1070_33_n_69, sub_1070_33_n_70, sub_1070_33_n_71,
     sub_1070_33_n_72, sub_1070_33_n_73, sub_1070_33_n_74, sub_1070_33_n_75,
     sub_1070_33_n_76, sub_1070_33_n_77, sub_1070_33_n_78, sub_1070_33_n_79,
     sub_1070_33_n_80, sub_1070_33_n_81, sub_1070_33_n_82, sub_1070_33_n_83,
     sub_1070_33_n_84, sub_1070_33_n_85, sub_1070_33_n_86, sub_1070_33_n_87,
     sub_1070_33_n_88, sub_1070_33_n_89, sub_1070_33_n_90, sub_1070_33_n_91,
     sub_1070_33_n_92, sub_1070_33_n_93, sub_1070_33_n_94, sub_1070_33_n_95,
     sub_1070_33_n_96, sub_1070_33_n_97, sub_1070_33_n_98, sub_1070_33_n_99,
     sub_1070_33_n_100, sub_1070_33_n_101, sub_1070_33_n_102, sub_1070_33_n_103,
     sub_1070_33_n_104, sub_1070_33_n_105, sub_1070_33_n_106, sub_1070_33_n_107,
     sub_1070_33_n_108, sub_1070_33_n_110, sub_1070_33_n_111, sub_1070_33_n_112,
     sub_1070_33_n_113, sub_1070_33_n_114, sub_1070_33_n_115, sub_1070_33_n_116,
     sub_1070_33_n_117, sub_1070_33_n_118, sub_1070_33_n_119, sub_1070_33_n_120,
     sub_1070_33_n_121, sub_1070_33_n_122, sub_1070_33_n_123, sub_1070_33_n_124,
     sub_1070_33_n_125, sub_1070_33_n_126, sub_1070_33_n_127, sub_1070_33_n_128,
     sub_1070_33_n_129, sub_1070_33_n_130, sub_1070_33_n_131, sub_1070_33_n_132,
     sub_1070_33_n_133, sub_1070_33_n_134, sub_1070_33_n_135, sub_1070_33_n_136,
     sub_1070_33_n_137, sub_1070_33_n_138, sub_1070_33_n_139, sub_1070_33_n_140,
     sub_1070_33_n_141, sub_1070_33_n_142, sub_1070_33_n_143, sub_1070_33_n_144,
     sub_1070_33_n_145, sub_1070_33_n_146, sub_1070_33_n_147, sub_1070_33_n_148,
     sub_1070_33_n_149, sub_1070_33_n_150, sub_1070_33_n_151, sub_1070_33_n_152,
     sub_1070_33_n_153, sub_1070_33_n_154, sub_1070_33_n_155, sub_1070_33_n_156,
     sub_1070_33_n_157, sub_1070_33_n_158, sub_1070_33_n_159, sub_1070_33_n_160,
     sub_1070_33_n_161, sub_1070_33_n_162, sub_1070_33_n_163, sub_1070_33_n_164,
     sub_1070_33_n_165, sub_1070_33_n_166, sub_1070_33_n_167, sub_1070_33_n_168,
     sub_1070_33_n_169, sub_1070_33_n_170, sub_1070_33_n_172, sub_1070_33_n_173,
     sub_1070_33_n_174, sub_1070_33_n_175, sub_1070_33_n_176, sub_1070_33_n_177,
     sub_1070_33_n_178, sub_1070_33_n_179, sub_1070_33_n_180, sub_1070_33_n_181,
     sub_1070_33_n_182, sub_1070_33_n_183, sub_1070_33_n_184, sub_1070_33_n_185,
     sub_1070_33_n_186, sub_1070_33_n_188, sub_1070_33_n_189, sub_1070_33_n_190,
     sub_1070_33_n_191, sub_1070_33_n_192, sub_1070_33_n_195, sub_1070_33_n_196,
     sub_1070_33_n_197, sub_1070_33_n_198, sub_1070_33_n_199, sub_1070_33_n_200,
     sub_1070_33_n_201, sub_1070_33_n_202, sub_1070_33_n_206, sub_1070_33_n_207,
     sub_1070_33_n_208, sub_1070_33_n_209, sub_1070_33_n_210, sub_1070_33_n_211,
     sub_1070_33_n_212, sub_1070_33_n_213, sub_1070_33_n_214, sub_1070_33_n_220,
     sub_1070_33_n_221, sub_1070_33_n_222, sub_1070_33_n_223, sub_1070_33_n_224,
     sub_1070_33_n_225, sub_1070_33_n_236, sub_1070_33_n_237, sub_1070_33_n_238,
     sub_1100_32_n_0, sub_1100_32_n_1, sub_1100_32_n_2, sub_1100_32_n_3,
     sub_1100_32_n_4, sub_1100_32_n_5, sub_1100_32_n_6, sub_1100_32_n_7,
     sub_1100_32_n_8, sub_1100_32_n_9, sub_1100_32_n_10, sub_1100_32_n_11,
     sub_1100_32_n_12, sub_1100_32_n_13, sub_1100_32_n_14, sub_1100_32_n_15,
     sub_1100_32_n_16, sub_1100_32_n_17, sub_1100_32_n_18, sub_1100_32_n_19,
     sub_1100_32_n_20, sub_1100_32_n_21, sub_1100_32_n_22, sub_1100_32_n_23,
     sub_1100_32_n_24, sub_1100_32_n_25, sub_1100_32_n_26, sub_1100_32_n_27,
     sub_1100_32_n_28, sub_1100_32_n_29, sub_1100_32_n_30, sub_1100_32_n_31,
     sub_1100_32_n_32, sub_1100_32_n_33, sub_1100_32_n_34, sub_1100_32_n_35,
     sub_1100_32_n_36, sub_1100_32_n_37, sub_1100_32_n_38, sub_1100_32_n_39,
     sub_1100_32_n_40, sub_1100_32_n_41, sub_1100_32_n_42, sub_1100_32_n_43,
     sub_1100_32_n_44, sub_1100_32_n_46, sub_1100_32_n_47, sub_1100_32_n_48,
     sub_1100_32_n_49, sub_1100_32_n_50, sub_1100_32_n_51, sub_1100_32_n_52,
     sub_1100_32_n_53, sub_1100_32_n_54, sub_1100_32_n_55, sub_1100_32_n_56,
     sub_1100_32_n_57, sub_1100_32_n_58, sub_1100_32_n_59, sub_1100_32_n_60,
     sub_1100_32_n_61, sub_1100_32_n_62, sub_1100_32_n_63, sub_1100_32_n_64,
     sub_1100_32_n_65, sub_1100_32_n_66, sub_1100_32_n_67, sub_1100_32_n_68,
     sub_1100_32_n_69, sub_1100_32_n_70, sub_1100_32_n_71, sub_1100_32_n_72,
     sub_1100_32_n_73, sub_1100_32_n_74, sub_1100_32_n_75, sub_1100_32_n_76,
     sub_1100_32_n_77, sub_1100_32_n_78, sub_1100_32_n_79, sub_1100_32_n_80,
     sub_1100_32_n_81, sub_1100_32_n_82, sub_1100_32_n_83, sub_1100_32_n_84,
     sub_1100_32_n_85, sub_1100_32_n_86, sub_1100_32_n_87, sub_1100_32_n_88,
     sub_1100_32_n_89, sub_1100_32_n_90, sub_1100_32_n_91, sub_1100_32_n_92,
     sub_1100_32_n_93, sub_1100_32_n_94, sub_1100_32_n_95, sub_1100_32_n_96,
     sub_1100_32_n_97, sub_1100_32_n_98, sub_1100_32_n_99, sub_1100_32_n_100,
     sub_1100_32_n_101, sub_1100_32_n_102, sub_1100_32_n_103, sub_1100_32_n_104,
     sub_1100_32_n_105, sub_1100_32_n_106, sub_1100_32_n_107, sub_1100_32_n_108,
     sub_1100_32_n_109, sub_1100_32_n_110, sub_1100_32_n_111, sub_1100_32_n_112,
     sub_1100_32_n_113, sub_1100_32_n_114, sub_1100_32_n_115, sub_1100_32_n_116,
     sub_1100_32_n_117, sub_1100_32_n_118, sub_1100_32_n_119, sub_1100_32_n_120,
     sub_1100_32_n_121, sub_1100_32_n_122, sub_1100_32_n_123, sub_1100_32_n_124,
     sub_1100_32_n_125, sub_1100_32_n_126, sub_1100_32_n_128, sub_1100_32_n_129,
     sub_1100_32_n_130, sub_1100_32_n_131, sub_1100_32_n_132, sub_1100_32_n_133,
     sub_1100_32_n_134, sub_1100_32_n_135, sub_1100_32_n_136, sub_1100_32_n_137,
     sub_1100_32_n_138, sub_1100_32_n_139, sub_1100_32_n_140, sub_1100_32_n_141,
     sub_1100_32_n_142, sub_1100_32_n_143, sub_1100_32_n_144, sub_1100_32_n_145,
     sub_1100_32_n_146, sub_1100_32_n_147, sub_1100_32_n_148, sub_1100_32_n_149,
     sub_1100_32_n_150, sub_1100_32_n_151, sub_1100_32_n_152, sub_1100_32_n_153,
     sub_1100_32_n_154, sub_1100_32_n_155, sub_1100_32_n_156, sub_1100_32_n_157,
     sub_1100_32_n_158, sub_1100_32_n_159, sub_1100_32_n_160, sub_1100_32_n_161,
     sub_1100_32_n_162, sub_1100_32_n_163, sub_1100_32_n_164, sub_1100_32_n_165,
     sub_1100_32_n_166, sub_1100_32_n_167, sub_1100_32_n_168, sub_1100_32_n_169,
     sub_1100_32_n_170, sub_1100_32_n_171, sub_1100_32_n_172, sub_1100_32_n_173,
     sub_1100_32_n_174, sub_1100_32_n_175, sub_1100_32_n_176, sub_1100_32_n_177,
     sub_1100_32_n_178, sub_1100_32_n_179, sub_1100_32_n_180, sub_1100_32_n_181,
     sub_1100_32_n_182, sub_1100_32_n_183, sub_1100_32_n_184, sub_1100_32_n_185,
     sub_1100_32_n_186, sub_1100_32_n_187, sub_1100_32_n_188, sub_1100_32_n_189,
     sub_1100_32_n_190, sub_1100_32_n_191, sub_1100_32_n_192, sub_1100_32_n_193,
     sub_1100_32_n_194, sub_1100_32_n_195, sub_1100_32_n_196, sub_1100_32_n_197,
     sub_1100_32_n_198, sub_1100_32_n_200, sub_1100_32_n_201, sub_1100_32_n_202,
     sub_1100_32_n_203, sub_1100_32_n_205, sub_1100_32_n_206, sub_1100_32_n_207,
     sub_1100_32_n_208, sub_1100_32_n_209, sub_1100_32_n_212, sub_1100_32_n_213,
     sub_1100_32_n_214, sub_1100_32_n_215, sub_1100_32_n_219, sub_1100_32_n_220,
     sub_1100_32_n_221, sub_1100_32_n_222, sub_1100_32_n_223, sub_1100_32_n_224,
     sub_1100_32_n_225, sub_1100_32_n_226, sub_1100_32_n_227, sub_1100_32_n_228,
     sub_1100_32_n_234, sub_1100_32_n_235, sub_1100_32_n_236, sub_1100_32_n_237,
     sub_1100_32_n_238, sub_1100_32_n_239, sub_1100_32_n_248, sub_1100_32_n_249,
     sub_1100_32_n_250, sub_1100_32_n_251, sub_1100_32_n_252, sub_1100_32_n_260,
     sub_1100_32_n_261, sub_1100_32_n_262, sub_1130_31_n_0, sub_1130_31_n_1,
     sub_1130_31_n_2, sub_1130_31_n_3, sub_1130_31_n_4, sub_1130_31_n_5,
     sub_1130_31_n_6, sub_1130_31_n_7, sub_1130_31_n_8, sub_1130_31_n_9,
     sub_1130_31_n_10, sub_1130_31_n_11, sub_1130_31_n_12, sub_1130_31_n_13,
     sub_1130_31_n_14, sub_1130_31_n_15, sub_1130_31_n_16, sub_1130_31_n_17,
     sub_1130_31_n_18, sub_1130_31_n_19, sub_1130_31_n_20, sub_1130_31_n_21,
     sub_1130_31_n_22, sub_1130_31_n_23, sub_1130_31_n_24, sub_1130_31_n_25,
     sub_1130_31_n_26, sub_1130_31_n_27, sub_1130_31_n_28, sub_1130_31_n_29,
     sub_1130_31_n_30, sub_1130_31_n_31, sub_1130_31_n_32, sub_1130_31_n_33,
     sub_1130_31_n_34, sub_1130_31_n_35, sub_1130_31_n_36, sub_1130_31_n_37,
     sub_1130_31_n_38, sub_1130_31_n_39, sub_1130_31_n_40, sub_1130_31_n_41,
     sub_1130_31_n_42, sub_1130_31_n_43, sub_1130_31_n_44, sub_1130_31_n_45,
     sub_1130_31_n_46, sub_1130_31_n_47, sub_1130_31_n_48, sub_1130_31_n_49,
     sub_1130_31_n_50, sub_1130_31_n_51, sub_1130_31_n_52, sub_1130_31_n_53,
     sub_1130_31_n_54, sub_1130_31_n_55, sub_1130_31_n_56, sub_1130_31_n_57,
     sub_1130_31_n_58, sub_1130_31_n_59, sub_1130_31_n_60, sub_1130_31_n_61,
     sub_1130_31_n_62, sub_1130_31_n_63, sub_1130_31_n_64, sub_1130_31_n_65,
     sub_1130_31_n_66, sub_1130_31_n_67, sub_1130_31_n_68, sub_1130_31_n_69,
     sub_1130_31_n_70, sub_1130_31_n_71, sub_1130_31_n_72, sub_1130_31_n_73,
     sub_1130_31_n_74, sub_1130_31_n_75, sub_1130_31_n_76, sub_1130_31_n_77,
     sub_1130_31_n_78, sub_1130_31_n_79, sub_1130_31_n_80, sub_1130_31_n_81,
     sub_1130_31_n_82, sub_1130_31_n_83, sub_1130_31_n_84, sub_1130_31_n_85,
     sub_1130_31_n_86, sub_1130_31_n_87, sub_1130_31_n_88, sub_1130_31_n_89,
     sub_1130_31_n_90, sub_1130_31_n_91, sub_1130_31_n_92, sub_1130_31_n_93,
     sub_1130_31_n_94, sub_1130_31_n_95, sub_1130_31_n_96, sub_1130_31_n_97,
     sub_1130_31_n_98, sub_1130_31_n_99, sub_1130_31_n_100, sub_1130_31_n_101,
     sub_1130_31_n_102, sub_1130_31_n_103, sub_1130_31_n_104, sub_1130_31_n_105,
     sub_1130_31_n_106, sub_1130_31_n_107, sub_1130_31_n_108, sub_1130_31_n_110,
     sub_1130_31_n_111, sub_1130_31_n_112, sub_1130_31_n_113, sub_1130_31_n_114,
     sub_1130_31_n_115, sub_1130_31_n_116, sub_1130_31_n_117, sub_1130_31_n_118,
     sub_1130_31_n_119, sub_1130_31_n_120, sub_1130_31_n_121, sub_1130_31_n_122,
     sub_1130_31_n_123, sub_1130_31_n_124, sub_1130_31_n_125, sub_1130_31_n_126,
     sub_1130_31_n_127, sub_1130_31_n_128, sub_1130_31_n_129, sub_1130_31_n_130,
     sub_1130_31_n_131, sub_1130_31_n_132, sub_1130_31_n_133, sub_1130_31_n_134,
     sub_1130_31_n_135, sub_1130_31_n_136, sub_1130_31_n_137, sub_1130_31_n_138,
     sub_1130_31_n_139, sub_1130_31_n_140, sub_1130_31_n_141, sub_1130_31_n_142,
     sub_1130_31_n_143, sub_1130_31_n_144, sub_1130_31_n_145, sub_1130_31_n_146,
     sub_1130_31_n_147, sub_1130_31_n_148, sub_1130_31_n_149, sub_1130_31_n_150,
     sub_1130_31_n_151, sub_1130_31_n_152, sub_1130_31_n_153, sub_1130_31_n_154,
     sub_1130_31_n_155, sub_1130_31_n_156, sub_1130_31_n_157, sub_1130_31_n_158,
     sub_1130_31_n_159, sub_1130_31_n_160, sub_1130_31_n_161, sub_1130_31_n_162,
     sub_1130_31_n_163, sub_1130_31_n_164, sub_1130_31_n_165, sub_1130_31_n_166,
     sub_1130_31_n_167, sub_1130_31_n_168, sub_1130_31_n_169, sub_1130_31_n_170,
     sub_1130_31_n_171, sub_1130_31_n_172, sub_1130_31_n_173, sub_1130_31_n_174,
     sub_1130_31_n_175, sub_1130_31_n_176, sub_1130_31_n_177, sub_1130_31_n_178,
     sub_1130_31_n_179, sub_1130_31_n_180, sub_1130_31_n_182, sub_1130_31_n_183,
     sub_1130_31_n_184, sub_1130_31_n_185, sub_1130_31_n_186, sub_1130_31_n_187,
     sub_1130_31_n_189, sub_1130_31_n_190, sub_1130_31_n_191, sub_1130_31_n_192,
     sub_1130_31_n_193, sub_1130_31_n_196, sub_1130_31_n_197, sub_1130_31_n_198,
     sub_1130_31_n_199, sub_1130_31_n_200, sub_1130_31_n_201, sub_1130_31_n_202,
     sub_1130_31_n_206, sub_1130_31_n_207, sub_1130_31_n_208, sub_1130_31_n_209,
     sub_1130_31_n_210, sub_1130_31_n_211, sub_1130_31_n_212, sub_1130_31_n_213,
     sub_1130_31_n_219, sub_1130_31_n_220, sub_1130_31_n_222, sub_1130_31_n_223,
     sub_1130_31_n_224, sub_1130_31_n_232, sub_1130_31_n_233, sub_1130_31_n_234,
     sub_1130_31_n_235, sub_1130_31_n_236, sub_1130_31_n_237, sub_1130_31_n_238,
     sub_1130_31_n_239, sub_1130_31_n_247, sub_1130_31_n_248, sub_1130_31_n_249,
     sub_1130_31_n_250, sub_1160_30_n_0, sub_1160_30_n_1, sub_1160_30_n_2,
     sub_1160_30_n_3, sub_1160_30_n_4, sub_1160_30_n_6, sub_1160_30_n_7,
     sub_1160_30_n_8, sub_1160_30_n_9, sub_1160_30_n_10, sub_1160_30_n_11,
     sub_1160_30_n_12, sub_1160_30_n_13, sub_1160_30_n_14, sub_1160_30_n_15,
     sub_1160_30_n_16, sub_1160_30_n_17, sub_1160_30_n_18, sub_1160_30_n_19,
     sub_1160_30_n_20, sub_1160_30_n_21, sub_1160_30_n_22, sub_1160_30_n_23,
     sub_1160_30_n_24, sub_1160_30_n_25, sub_1160_30_n_26, sub_1160_30_n_27,
     sub_1160_30_n_28, sub_1160_30_n_29, sub_1160_30_n_30, sub_1160_30_n_31,
     sub_1160_30_n_32, sub_1160_30_n_33, sub_1160_30_n_34, sub_1160_30_n_35,
     sub_1160_30_n_36, sub_1160_30_n_37, sub_1160_30_n_38, sub_1160_30_n_39,
     sub_1160_30_n_40, sub_1160_30_n_41, sub_1160_30_n_42, sub_1160_30_n_43,
     sub_1160_30_n_44, sub_1160_30_n_45, sub_1160_30_n_46, sub_1160_30_n_47,
     sub_1160_30_n_48, sub_1160_30_n_49, sub_1160_30_n_50, sub_1160_30_n_51,
     sub_1160_30_n_52, sub_1160_30_n_53, sub_1160_30_n_54, sub_1160_30_n_55,
     sub_1160_30_n_56, sub_1160_30_n_57, sub_1160_30_n_58, sub_1160_30_n_59,
     sub_1160_30_n_60, sub_1160_30_n_61, sub_1160_30_n_62, sub_1160_30_n_63,
     sub_1160_30_n_64, sub_1160_30_n_65, sub_1160_30_n_66, sub_1160_30_n_67,
     sub_1160_30_n_68, sub_1160_30_n_69, sub_1160_30_n_70, sub_1160_30_n_71,
     sub_1160_30_n_72, sub_1160_30_n_73, sub_1160_30_n_74, sub_1160_30_n_75,
     sub_1160_30_n_76, sub_1160_30_n_77, sub_1160_30_n_78, sub_1160_30_n_79,
     sub_1160_30_n_80, sub_1160_30_n_81, sub_1160_30_n_82, sub_1160_30_n_83,
     sub_1160_30_n_84, sub_1160_30_n_85, sub_1160_30_n_86, sub_1160_30_n_87,
     sub_1160_30_n_88, sub_1160_30_n_89, sub_1160_30_n_90, sub_1160_30_n_91,
     sub_1160_30_n_92, sub_1160_30_n_93, sub_1160_30_n_94, sub_1160_30_n_95,
     sub_1160_30_n_96, sub_1160_30_n_97, sub_1160_30_n_98, sub_1160_30_n_99,
     sub_1160_30_n_100, sub_1160_30_n_101, sub_1160_30_n_102, sub_1160_30_n_103,
     sub_1160_30_n_104, sub_1160_30_n_105, sub_1160_30_n_106, sub_1160_30_n_107,
     sub_1160_30_n_108, sub_1160_30_n_109, sub_1160_30_n_110, sub_1160_30_n_111,
     sub_1160_30_n_112, sub_1160_30_n_113, sub_1160_30_n_114, sub_1160_30_n_115,
     sub_1160_30_n_116, sub_1160_30_n_117, sub_1160_30_n_118, sub_1160_30_n_119,
     sub_1160_30_n_120, sub_1160_30_n_121, sub_1160_30_n_122, sub_1160_30_n_123,
     sub_1160_30_n_124, sub_1160_30_n_125, stall, clk, n_756, n_757, n_758,
     n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769,
     n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780,
     n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_829, n_830, n_831, n_832,
     n_833, n_834, n_835, n_836, n_838, n_839, n_840, n_841, n_842, n_843, n_844,
     n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855,
     n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866,
     n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877,
     n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_889,
     n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900,
     n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911,
     n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922,
     n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933,
     n_934, n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944,
     n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955,
     n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966,
     n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977,
     n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988,
     n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999,
     n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008,
     n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017,
     n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026,
     n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035,
     n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044,
     n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053,
     n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062,
     n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071,
     n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080,
     n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089,
     n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098,
     n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107,
     n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116,
     n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125,
     n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134,
     n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143,
     n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152,
     n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161,
     n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170,
     n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179,
     n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188,
     n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197,
     n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206,
     n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215,
     n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224,
     n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233,
     n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242,
     n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251,
     n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260,
     n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269,
     n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278,
     n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287,
     n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296,
     n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305,
     n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314,
     n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323,
     n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332,
     n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341,
     n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350,
     n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359,
     n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368,
     n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377,
     n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, clr, Q_0_, Q_1_, Q_2_, Q_3_,
     Q_4_, Q_5_, Q_6_, Q_7_, R_1_0_, R_1_1_, R_1_2_, R_1_3_, R_1_4_, R_1_5_,
     R_1_6_, R_1_7_, R_1_8_, R_1_9_, R_1_10_, R_1_11_, R_1_12_, R_1_13_, R_1_14_,
     R_1_15_, R_1_16_, R_1_17_, R_1_18_, R_1_19_, R_1_20_, R_1_21_, R_1_22_,
     R_1_23_, R_1_24_, R_1_25_, R_1_26_, R_1_27_, R_1_28_, R_1_29_, R_1_30_,
     R_2_0_, R_2_1_, R_2_2_, R_2_3_, R_2_4_, R_2_5_, R_2_6_, R_2_7_, R_2_8_,
     R_2_9_, R_2_10_, R_2_11_, R_2_12_, R_2_13_, R_2_14_, R_2_15_, R_2_16_,
     R_2_17_, R_2_18_, R_2_19_, R_2_20_, R_2_21_, R_2_22_, R_2_23_, R_2_24_,
     R_2_25_, R_2_26_, R_2_27_, R_2_28_, R_2_29_, R_3_0_, R_3_1_, R_3_2_, R_3_3_,
     R_3_4_, R_3_5_, R_3_6_, R_3_7_, R_3_8_, R_3_9_, R_3_10_, R_3_11_, R_3_12_,
     R_3_13_, R_3_14_, R_3_15_, R_3_16_, R_3_17_, R_3_18_, R_3_19_, R_3_20_,
     R_3_21_, R_3_22_, R_3_23_, R_3_24_, R_3_25_, R_3_26_, R_3_27_, R_3_28_,
     R_4_0_, R_4_1_, R_4_2_, R_4_3_, R_4_4_, R_4_5_, R_4_6_, R_4_7_, R_4_8_,
     R_4_9_, R_4_10_, R_4_11_, R_4_12_, R_4_13_, R_4_14_, R_4_15_, R_4_16_,
     R_4_17_, R_4_18_, R_4_19_, R_4_20_, R_4_21_, R_4_22_, R_4_23_, R_4_24_,
     R_4_25_, R_4_26_, R_4_27_, R_5_0_, R_5_1_, R_5_2_, R_5_3_, R_5_4_, R_5_5_,
     R_5_6_, R_5_7_, R_5_8_, R_5_9_, R_5_10_, R_5_11_, R_5_12_, R_5_13_, R_5_14_,
     R_5_15_, R_5_16_, R_5_17_, R_5_18_, R_5_19_, R_5_20_, R_5_21_, R_5_22_,
     R_5_23_, R_5_24_, R_5_25_, R_5_26_, R_6_0_, R_6_1_, R_6_2_, R_6_3_, R_6_4_,
     R_6_5_, R_6_6_, R_6_7_, R_6_8_, R_6_9_, R_6_10_, R_6_11_, R_6_12_, R_6_13_,
     R_6_14_, R_6_15_, R_6_16_, R_6_17_, R_6_18_, R_6_19_, R_6_20_, R_6_21_,
     R_6_22_, R_6_23_, R_6_24_, R_6_25_, R_7_0_, R_7_1_, R_7_2_, R_7_3_, R_7_4_,
     R_7_5_, R_7_6_, R_7_7_, R_7_8_, R_7_9_, R_7_10_, R_7_11_, R_7_12_, R_7_13_,
     R_7_14_, R_7_15_, R_7_16_, R_7_17_, R_7_18_, R_7_19_, R_7_20_, R_7_21_,
     R_7_22_, R_7_23_, R_7_24_, R_8_0_, R_8_1_, R_8_2_, R_8_3_, R_8_4_, R_8_5_,
     R_8_6_, R_8_7_, R_8_8_, R_8_9_, R_8_10_, R_8_11_, R_8_12_, R_8_13_, R_8_14_,
     R_8_15_, R_8_16_, R_8_17_, R_8_18_, R_8_19_, R_8_20_, R_8_21_, R_8_22_,
     R_8_23_, R_9_0_, R_9_1_, R_9_2_, R_9_3_, R_9_4_, R_9_5_, R_9_6_, R_9_7_,
     R_9_8_, R_9_9_, R_9_10_, R_9_11_, R_9_12_, R_9_13_, R_9_14_, R_9_15_,
     R_9_16_, R_9_17_, R_9_18_, R_9_19_, R_9_20_, R_9_21_, R_9_22_, R_10_0_,
     R_10_1_, R_10_2_, R_10_3_, R_10_4_, R_10_5_, R_10_6_, R_10_7_, R_10_8_,
     R_10_9_, R_10_10_, R_10_11_, R_10_12_, R_10_13_, R_10_14_, R_10_15_,
     R_10_16_, R_10_17_, R_10_18_, R_10_19_, R_10_20_, R_10_21_, R_11_0_,
     R_11_1_, R_11_2_, R_11_3_, R_11_4_, R_11_5_, R_11_6_, R_11_7_, R_11_8_,
     R_11_9_, R_11_10_, R_11_11_, R_11_12_, R_11_13_, R_11_14_, R_11_15_,
     R_11_16_, R_11_17_, R_11_18_, R_11_19_, R_11_20_, R_12_0_, R_12_1_, R_12_2_,
     R_12_3_, R_12_4_, R_12_5_, R_12_6_, R_12_7_, R_12_8_, R_12_9_, R_12_10_,
     R_12_11_, R_12_12_, R_12_13_, R_12_14_, R_12_15_, R_12_16_, R_12_17_,
     R_12_18_, R_12_19_, R_13_0_, R_13_1_, R_13_2_, R_13_3_, R_13_4_, R_13_5_,
     R_13_6_, R_13_7_, R_13_8_, R_13_9_, R_13_10_, R_13_11_, R_13_12_, R_13_13_,
     R_13_14_, R_13_15_, R_13_16_, R_13_17_, R_13_18_, R_14_0_, R_14_1_, R_14_2_,
     R_14_3_, R_14_4_, R_14_5_, R_14_6_, R_14_7_, R_14_8_, R_14_9_, R_14_10_,
     R_14_11_, R_14_12_, R_14_13_, R_14_14_, R_14_15_, R_14_16_, R_14_17_,
     R_15_0_, R_15_1_, R_15_2_, R_15_3_, R_15_4_, R_15_5_, R_15_6_, R_15_7_,
     R_15_8_, R_15_9_, R_15_10_, R_15_11_, R_15_12_, R_15_13_, R_15_14_,
     R_15_15_, R_15_16_, R_16_0_, R_16_1_, R_16_2_, R_16_3_, R_16_4_, R_16_5_,
     R_16_6_, R_16_7_, R_16_8_, R_16_9_, R_16_10_, R_16_11_, R_16_12_, R_16_13_,
     R_16_14_, R_16_15_, R_17_0_, R_17_1_, R_17_2_, R_17_3_, R_17_4_, R_17_5_,
     R_17_6_, R_17_7_, R_17_8_, R_17_9_, R_17_10_, R_17_11_, R_17_12_, R_17_13_,
     R_17_14_, R_18_0_, R_18_1_, R_18_2_, R_18_3_, R_18_4_, R_18_5_, R_18_6_,
     R_18_7_, R_18_8_, R_18_9_, R_18_10_, R_18_11_, R_18_12_, R_18_13_, R_19_0_,
     R_19_1_, R_19_2_, R_19_3_, R_19_4_, R_19_5_, R_19_6_, R_19_7_, R_19_8_,
     R_19_9_, R_19_10_, R_19_11_, R_19_12_, R_20_0_, R_20_1_, R_20_2_, R_20_3_,
     R_20_4_, R_20_5_, R_20_6_, R_20_7_, R_20_8_, R_20_9_, R_20_10_, R_20_11_,
     R_21_0_, R_21_1_, R_21_2_, R_21_3_, R_21_4_, R_21_5_, R_21_6_, R_21_7_,
     R_21_8_, R_21_9_, R_21_10_, R_22_0_, R_22_1_, R_22_2_, R_22_3_, R_22_4_,
     R_22_5_, R_22_6_, R_22_7_, R_22_8_, R_22_9_, R_23_0_, R_23_1_, R_23_2_,
     R_23_3_, R_23_4_, R_23_5_, R_23_6_, R_23_7_, R_23_8_, R_24_0_, R_24_1_,
     R_24_2_, R_24_3_, R_24_4_, R_24_5_, R_24_6_, R_24_7_, R_25_0_, R_25_1_,
     R_25_2_, R_25_3_, R_25_4_, R_25_5_, R_25_6_, R_26_0_, R_26_1_, R_26_2_,
     R_26_3_, R_26_4_, R_26_5_, R_27_0_, R_27_1_, R_27_2_, R_27_3_, R_27_4_,
     R_28_0_, R_28_1_, R_28_2_, R_28_3_, R_29_0_, R_29_1_, R_29_2_, R_30_0_,
     R_30_1_, R_31_0_, T_0_32_, T_1_0_, T_1_1_, T_1_2_, T_1_3_, T_1_4_, T_1_5_,
     T_1_6_, T_1_7_, T_1_8_, T_1_9_, T_1_10_, T_1_11_, T_1_12_, T_1_13_, T_1_14_,
     T_1_15_, T_1_16_, T_1_17_, T_1_18_, T_1_19_, T_1_20_, T_1_21_, T_1_22_,
     T_1_23_, T_1_24_, T_1_25_, T_1_26_, T_1_27_, T_1_28_, T_1_29_, T_1_30_,
     T_1_32_, T_2_0_, T_2_1_, T_2_2_, T_2_3_, T_2_4_, T_2_5_, T_2_6_, T_2_7_,
     T_2_8_, T_2_9_, T_2_10_, T_2_11_, T_2_12_, T_2_13_, T_2_14_, T_2_15_,
     T_2_16_, T_2_17_, T_2_18_, T_2_19_, T_2_20_, T_2_21_, T_2_22_, T_2_23_,
     T_2_24_, T_2_25_, T_2_26_, T_2_27_, T_2_28_, T_2_29_, T_2_32_, T_3_0_,
     T_3_1_, T_3_2_, T_3_3_, T_3_4_, T_3_5_, T_3_6_, T_3_7_, T_3_8_, T_3_9_,
     T_3_10_, T_3_11_, T_3_12_, T_3_13_, T_3_14_, T_3_15_, T_3_16_, T_3_17_,
     T_3_18_, T_3_19_, T_3_20_, T_3_21_, T_3_22_, T_3_23_, T_3_24_, T_3_25_,
     T_3_26_, T_3_27_, T_3_28_, T_3_32_, T_4_0_, T_4_1_, T_4_2_, T_4_3_, T_4_4_,
     T_4_5_, T_4_6_, T_4_7_, T_4_8_, T_4_9_, T_4_10_, T_4_11_, T_4_12_, T_4_13_,
     T_4_14_, T_4_15_, T_4_16_, T_4_17_, T_4_18_, T_4_19_, T_4_20_, T_4_21_,
     T_4_22_, T_4_23_, T_4_24_, T_4_25_, T_4_26_, T_4_27_, T_4_32_, T_5_0_,
     T_5_1_, T_5_2_, T_5_3_, T_5_4_, T_5_5_, T_5_6_, T_5_7_, T_5_8_, T_5_9_,
     T_5_10_, T_5_11_, T_5_12_, T_5_13_, T_5_14_, T_5_15_, T_5_16_, T_5_17_,
     T_5_18_, T_5_19_, T_5_20_, T_5_21_, T_5_22_, T_5_23_, T_5_24_, T_5_25_,
     T_5_26_, T_5_32_, T_6_0_, T_6_1_, T_6_2_, T_6_3_, T_6_4_, T_6_5_, T_6_6_,
     T_6_7_, T_6_8_, T_6_9_, T_6_10_, T_6_11_, T_6_12_, T_6_13_, T_6_14_,
     T_6_15_, T_6_16_, T_6_17_, T_6_18_, T_6_19_, T_6_20_, T_6_21_, T_6_22_,
     T_6_23_, T_6_24_, T_6_25_, T_6_32_, T_7_0_, T_7_1_, T_7_2_, T_7_3_, T_7_4_,
     T_7_5_, T_7_6_, T_7_7_, T_7_8_, T_7_9_, T_7_10_, T_7_11_, T_7_12_, T_7_13_,
     T_7_14_, T_7_15_, T_7_16_, T_7_17_, T_7_18_, T_7_19_, T_7_20_, T_7_21_,
     T_7_22_, T_7_23_, T_7_24_, T_7_32_, T_8_0_, T_8_1_, T_8_2_, T_8_3_, T_8_4_,
     T_8_5_, T_8_6_, T_8_7_, T_8_8_, T_8_9_, T_8_10_, T_8_11_, T_8_12_, T_8_13_,
     T_8_14_, T_8_15_, T_8_16_, T_8_17_, T_8_18_, T_8_19_, T_8_20_, T_8_21_,
     T_8_22_, T_8_23_, T_8_32_, T_9_0_, T_9_1_, T_9_2_, T_9_3_, T_9_4_, T_9_5_,
     T_9_6_, T_9_7_, T_9_8_, T_9_9_, T_9_10_, T_9_11_, T_9_12_, T_9_13_, T_9_14_,
     T_9_15_, T_9_16_, T_9_17_, T_9_18_, T_9_19_, T_9_20_, T_9_21_, T_9_22_,
     T_9_32_, T_10_0_, T_10_1_, T_10_2_, T_10_3_, T_10_4_, T_10_5_, T_10_6_,
     T_10_7_, T_10_8_, T_10_9_, T_10_10_, T_10_11_, T_10_12_, T_10_13_, T_10_14_,
     T_10_15_, T_10_16_, T_10_17_, T_10_18_, T_10_19_, T_10_20_, T_10_21_,
     T_10_32_, T_11_0_, T_11_1_, T_11_2_, T_11_3_, T_11_4_, T_11_5_, T_11_6_,
     T_11_7_, T_11_8_, T_11_9_, T_11_10_, T_11_11_, T_11_12_, T_11_13_, T_11_14_,
     T_11_15_, T_11_16_, T_11_17_, T_11_18_, T_11_19_, T_11_20_, T_11_32_,
     T_12_0_, T_12_1_, T_12_2_, T_12_3_, T_12_4_, T_12_5_, T_12_6_, T_12_7_,
     T_12_8_, T_12_9_, T_12_10_, T_12_11_, T_12_12_, T_12_13_, T_12_14_,
     T_12_15_, T_12_16_, T_12_17_, T_12_18_, T_12_19_, T_12_32_, T_13_0_,
     T_13_1_, T_13_2_, T_13_3_, T_13_4_, T_13_5_, T_13_6_, T_13_7_, T_13_8_,
     T_13_9_, T_13_10_, T_13_11_, T_13_12_, T_13_13_, T_13_14_, T_13_15_,
     T_13_16_, T_13_17_, T_13_18_, T_13_32_, T_14_0_, T_14_1_, T_14_2_, T_14_3_,
     T_14_4_, T_14_5_, T_14_6_, T_14_7_, T_14_8_, T_14_9_, T_14_10_, T_14_11_,
     T_14_12_, T_14_13_, T_14_14_, T_14_15_, T_14_16_, T_14_17_, T_14_32_,
     T_15_0_, T_15_1_, T_15_2_, T_15_3_, T_15_4_, T_15_5_, T_15_6_, T_15_7_,
     T_15_8_, T_15_9_, T_15_10_, T_15_11_, T_15_12_, T_15_13_, T_15_14_,
     T_15_15_, T_15_16_, T_15_32_, T_16_0_, T_16_1_, T_16_2_, T_16_3_, T_16_4_,
     T_16_5_, T_16_6_, T_16_7_, T_16_8_, T_16_9_, T_16_10_, T_16_11_, T_16_12_,
     T_16_13_, T_16_14_, T_16_15_, T_16_32_, T_17_0_, T_17_1_, T_17_2_, T_17_3_,
     T_17_4_, T_17_5_, T_17_6_, T_17_7_, T_17_8_, T_17_9_, T_17_10_, T_17_11_,
     T_17_12_, T_17_13_, T_17_14_, T_17_32_, T_18_0_, T_18_1_, T_18_2_, T_18_3_,
     T_18_4_, T_18_5_, T_18_6_, T_18_7_, T_18_8_, T_18_9_, T_18_10_, T_18_11_,
     T_18_12_, T_18_13_, T_18_32_, T_19_0_, T_19_1_, T_19_2_, T_19_3_, T_19_4_,
     T_19_5_, T_19_6_, T_19_7_, T_19_8_, T_19_9_, T_19_10_, T_19_11_, T_19_12_,
     T_19_32_, T_20_0_, T_20_1_, T_20_2_, T_20_3_, T_20_4_, T_20_5_, T_20_6_,
     T_20_7_, T_20_8_, T_20_9_, T_20_10_, T_20_11_, T_20_32_, T_21_0_, T_21_1_,
     T_21_2_, T_21_3_, T_21_4_, T_21_5_, T_21_6_, T_21_7_, T_21_8_, T_21_9_,
     T_21_10_, T_21_32_, T_22_0_, T_22_1_, T_22_2_, T_22_3_, T_22_4_, T_22_5_,
     T_22_6_, T_22_7_, T_22_8_, T_22_9_, T_22_32_, T_23_0_, T_23_1_, T_23_2_,
     T_23_3_, T_23_4_, T_23_5_, T_23_6_, T_23_7_, T_23_8_, T_23_32_, T_24_0_,
     T_24_1_, T_24_2_, T_24_3_, T_24_4_, T_24_5_, T_24_6_, T_24_7_, T_24_32_,
     T_25_0_, T_25_1_, T_25_2_, T_25_3_, T_25_4_, T_25_5_, T_25_6_, T_25_32_,
     T_26_0_, T_26_1_, T_26_2_, T_26_3_, T_26_4_, T_26_5_, T_26_32_, T_27_0_,
     T_27_1_, T_27_2_, T_27_3_, T_27_4_, T_27_32_, T_28_0_, T_28_1_, T_28_2_,
     T_28_3_, T_28_32_, T_29_0_, T_29_1_, T_29_2_, T_29_32_, T_30_0_, T_30_1_,
     T_30_32_, T_31_0_, T_31_32_;
assign n_756 = Q_7_;
assign n_757 = Q_6_;
assign n_758 = Q_5_;
assign n_759 = Q_4_;
assign n_760 = Q_3_;
assign n_761 = Q_2_;
assign n_762 = Q_1_;
assign n_763 = Q_0_;
assign n_764 = n_756;
assign n_765 = n_757;
assign n_766 = n_758;
assign n_767 = n_759;
assign n_768 = n_760;
assign n_769 = n_761;
assign n_770 = n_762;
assign n_771 = n_763;
assign n_772 = n_764;
assign n_773 = n_765;
assign n_774 = n_766;
assign n_775 = n_767;
assign n_776 = n_768;
assign n_777 = n_769;
assign n_778 = n_770;
assign n_779 = n_771;
assign n_780 = n_772;
assign n_781 = n_773;
assign n_782 = n_774;
assign n_783 = n_775;
assign n_784 = n_776;
assign n_785 = n_777;
assign n_786 = n_778;
assign n_787 = n_779;
assign {out1[5]} = n_782;
assign {out1[4]} = n_783;
assign {out1[3]} = n_784;
assign {out1[2]} = n_785;
assign {out1[1]} = n_786;
assign {out1[0]} = n_787;
reg cadence_register_n_829;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_829 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_829 <= in1[30];
    end
 end
 assign n_829 = cadence_register_n_829;
reg cadence_register_n_830;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_830 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_830 <= n_829;
    end
 end
 assign n_830 = cadence_register_n_830;
reg cadence_register_n_831;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_831 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_831 <= n_830;
    end
 end
 assign n_831 = cadence_register_n_831;
reg cadence_register_n_832;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_832 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_832 <= n_831;
    end
 end
 assign n_832 = cadence_register_n_832;
reg cadence_register_n_833;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_833 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_833 <= n_832;
    end
 end
 assign n_833 = cadence_register_n_833;
reg cadence_register_n_834;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_834 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_834 <= sub_1040_34_n_116;
    end
 end
 assign n_834 = cadence_register_n_834;
reg cadence_register_n_835;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_835 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_835 <= T_5_32_;
    end
 end
 assign n_835 = cadence_register_n_835;
reg cadence_register_n_836;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_836 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_836 <= R_5_1_;
    end
 end
 assign n_836 = cadence_register_n_836;
reg cadence_register_out1_7;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_out1_7 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_out1_7 <= n_780;
    end
 end
 assign out1[7] = cadence_register_out1_7;
reg cadence_register_n_838;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_838 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_838 <= R_5_9_;
    end
 end
 assign n_838 = cadence_register_n_838;
reg cadence_register_n_839;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_839 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_839 <= sub_1040_34_n_6;
    end
 end
 assign n_839 = cadence_register_n_839;
reg cadence_register_n_840;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_840 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_840 <= sub_1040_34_n_84;
    end
 end
 assign n_840 = cadence_register_n_840;
reg cadence_register_n_841;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_841 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_841 <= R_5_8_;
    end
 end
 assign n_841 = cadence_register_n_841;
reg cadence_register_n_842;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_842 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_842 <= R_5_14_;
    end
 end
 assign n_842 = cadence_register_n_842;
reg cadence_register_n_843;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_843 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_843 <= R_5_18_;
    end
 end
 assign n_843 = cadence_register_n_843;
reg cadence_register_n_844;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_844 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_844 <= sub_1040_34_n_44;
    end
 end
 assign n_844 = cadence_register_n_844;
reg cadence_register_n_845;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_845 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_845 <= sub_1040_34_n_97;
    end
 end
 assign n_845 = cadence_register_n_845;
reg cadence_register_n_846;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_846 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_846 <= R_5_17_;
    end
 end
 assign n_846 = cadence_register_n_846;
reg cadence_register_n_847;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_847 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_847 <= sub_1040_34_n_101;
    end
 end
 assign n_847 = cadence_register_n_847;
reg cadence_register_n_848;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_848 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_848 <= sub_1040_34_n_81;
    end
 end
 assign n_848 = cadence_register_n_848;
reg cadence_register_n_849;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_849 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_849 <= R_5_16_;
    end
 end
 assign n_849 = cadence_register_n_849;
reg cadence_register_n_850;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_850 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_850 <= sub_1040_34_n_69;
    end
 end
 assign n_850 = cadence_register_n_850;
reg cadence_register_n_851;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_851 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_851 <= sub_1040_34_n_9;
    end
 end
 assign n_851 = cadence_register_n_851;
reg cadence_register_n_852;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_852 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_852 <= sub_1040_34_n_68;
    end
 end
 assign n_852 = cadence_register_n_852;
reg cadence_register_n_853;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_853 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_853 <= R_5_15_;
    end
 end
 assign n_853 = cadence_register_n_853;
reg cadence_register_n_854;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_854 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_854 <= R_5_19_;
    end
 end
 assign n_854 = cadence_register_n_854;
reg cadence_register_n_855;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_855 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_855 <= R_5_24_;
    end
 end
 assign n_855 = cadence_register_n_855;
reg cadence_register_n_856;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_856 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_856 <= R_5_21_;
    end
 end
 assign n_856 = cadence_register_n_856;
reg cadence_register_n_857;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_857 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_857 <= sub_1040_34_n_71;
    end
 end
 assign n_857 = cadence_register_n_857;
reg cadence_register_n_858;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_858 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_858 <= sub_1040_34_n_65;
    end
 end
 assign n_858 = cadence_register_n_858;
reg cadence_register_n_859;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_859 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_859 <= sub_1040_34_n_47;
    end
 end
 assign n_859 = cadence_register_n_859;
reg cadence_register_n_860;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_860 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_860 <= sub_1040_34_n_49;
    end
 end
 assign n_860 = cadence_register_n_860;
reg cadence_register_n_861;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_861 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_861 <= R_5_12_;
    end
 end
 assign n_861 = cadence_register_n_861;
reg cadence_register_n_862;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_862 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_862 <= R_5_13_;
    end
 end
 assign n_862 = cadence_register_n_862;
reg cadence_register_n_863;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_863 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_863 <= sub_1040_34_n_2;
    end
 end
 assign n_863 = cadence_register_n_863;
reg cadence_register_n_864;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_864 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_864 <= sub_1040_34_n_106;
    end
 end
 assign n_864 = cadence_register_n_864;
reg cadence_register_n_865;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_865 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_865 <= sub_1040_34_n_95;
    end
 end
 assign n_865 = cadence_register_n_865;
reg cadence_register_n_866;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_866 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_866 <= sub_1040_34_n_83;
    end
 end
 assign n_866 = cadence_register_n_866;
reg cadence_register_n_867;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_867 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_867 <= R_5_22_;
    end
 end
 assign n_867 = cadence_register_n_867;
reg cadence_register_n_868;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_868 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_868 <= sub_1040_34_n_105;
    end
 end
 assign n_868 = cadence_register_n_868;
reg cadence_register_n_869;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_869 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_869 <= sub_1040_34_n_109;
    end
 end
 assign n_869 = cadence_register_n_869;
reg cadence_register_n_870;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_870 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_870 <= R_5_26_;
    end
 end
 assign n_870 = cadence_register_n_870;
reg cadence_register_n_871;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_871 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_871 <= R_5_23_;
    end
 end
 assign n_871 = cadence_register_n_871;
reg cadence_register_n_872;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_872 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_872 <= R_5_7_;
    end
 end
 assign n_872 = cadence_register_n_872;
reg cadence_register_n_873;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_873 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_873 <= R_5_20_;
    end
 end
 assign n_873 = cadence_register_n_873;
reg cadence_register_n_874;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_874 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_874 <= sub_1040_34_n_98;
    end
 end
 assign n_874 = cadence_register_n_874;
reg cadence_register_n_875;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_875 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_875 <= R_5_25_;
    end
 end
 assign n_875 = cadence_register_n_875;
reg cadence_register_n_876;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_876 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_876 <= sub_1040_34_n_23;
    end
 end
 assign n_876 = cadence_register_n_876;
reg cadence_register_n_877;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_877 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_877 <= sub_1040_34_n_48;
    end
 end
 assign n_877 = cadence_register_n_877;
reg cadence_register_n_878;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_878 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_878 <= sub_1040_34_n_17;
    end
 end
 assign n_878 = cadence_register_n_878;
reg cadence_register_n_879;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_879 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_879 <= R_5_5_;
    end
 end
 assign n_879 = cadence_register_n_879;
reg cadence_register_n_880;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_880 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_880 <= R_5_6_;
    end
 end
 assign n_880 = cadence_register_n_880;
reg cadence_register_n_881;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_881 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_881 <= sub_1040_34_n_110;
    end
 end
 assign n_881 = cadence_register_n_881;
reg cadence_register_n_882;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_882 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_882 <= sub_1040_34_n_8;
    end
 end
 assign n_882 = cadence_register_n_882;
reg cadence_register_n_883;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_883 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_883 <= R_5_4_;
    end
 end
 assign n_883 = cadence_register_n_883;
reg cadence_register_n_884;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_884 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_884 <= sub_1040_34_n_107;
    end
 end
 assign n_884 = cadence_register_n_884;
reg cadence_register_n_885;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_885 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_885 <= sub_1040_34_n_12;
    end
 end
 assign n_885 = cadence_register_n_885;
reg cadence_register_n_886;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_886 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_886 <= sub_1040_34_n_46;
    end
 end
 assign n_886 = cadence_register_n_886;
reg cadence_register_n_887;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_887 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_887 <= sub_1040_34_n_66;
    end
 end
 assign n_887 = cadence_register_n_887;
reg cadence_register_out1_6;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_out1_6 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_out1_6 <= n_781;
    end
 end
 assign out1[6] = cadence_register_out1_6;
reg cadence_register_n_889;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_889 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_889 <= R_5_11_;
    end
 end
 assign n_889 = cadence_register_n_889;
reg cadence_register_n_890;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_890 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_890 <= R_5_10_;
    end
 end
 assign n_890 = cadence_register_n_890;
reg cadence_register_n_891;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_891 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_891 <= sub_1040_34_n_7;
    end
 end
 assign n_891 = cadence_register_n_891;
reg cadence_register_n_892;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_892 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_892 <= sub_1040_34_n_96;
    end
 end
 assign n_892 = cadence_register_n_892;
reg cadence_register_n_893;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_893 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_893 <= sub_1040_34_n_70;
    end
 end
 assign n_893 = cadence_register_n_893;
reg cadence_register_n_894;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_894 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_894 <= R_5_2_;
    end
 end
 assign n_894 = cadence_register_n_894;
reg cadence_register_n_895;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_895 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_895 <= T_4_3_;
    end
 end
 assign n_895 = cadence_register_n_895;
reg cadence_register_n_896;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_896 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_896 <= sub_1040_34_n_75;
    end
 end
 assign n_896 = cadence_register_n_896;
reg cadence_register_n_897;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_897 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_897 <= sub_1040_34_n_183;
    end
 end
 assign n_897 = cadence_register_n_897;
reg cadence_register_n_898;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_898 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_898 <= R_5_3_;
    end
 end
 assign n_898 = cadence_register_n_898;
reg cadence_register_n_899;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_899 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_899 <= sub_1040_34_n_11;
    end
 end
 assign n_899 = cadence_register_n_899;
reg cadence_register_n_900;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_900 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_900 <= sub_1040_34_n_10;
    end
 end
 assign n_900 = cadence_register_n_900;
reg cadence_register_n_901;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_901 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_901 <= R_5_0_;
    end
 end
 assign n_901 = cadence_register_n_901;
reg cadence_register_n_902;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_902 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_902 <= T_4_1_;
    end
 end
 assign n_902 = cadence_register_n_902;
reg cadence_register_n_903;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_903 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_903 <= T_4_2_;
    end
 end
 assign n_903 = cadence_register_n_903;
reg cadence_register_n_904;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_904 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_904 <= sub_1040_34_n_151;
    end
 end
 assign n_904 = cadence_register_n_904;
reg cadence_register_n_905;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_905 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_905 <= sub_1040_34_n_16;
    end
 end
 assign n_905 = cadence_register_n_905;
reg cadence_register_n_906;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_906 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_906 <= sub_1040_34_n_18;
    end
 end
 assign n_906 = cadence_register_n_906;
reg cadence_register_n_907;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_907 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_907 <= R_10_17_;
    end
 end
 assign n_907 = cadence_register_n_907;
reg cadence_register_n_908;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_908 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_908 <= sub_890_40_n_42;
    end
 end
 assign n_908 = cadence_register_n_908;
reg cadence_register_n_909;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_909 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_909 <= sub_890_40_n_179;
    end
 end
 assign n_909 = cadence_register_n_909;
reg cadence_register_n_910;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_910 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_910 <= R_10_4_;
    end
 end
 assign n_910 = cadence_register_n_910;
reg cadence_register_n_911;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_911 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_911 <= T_9_7_;
    end
 end
 assign n_911 = cadence_register_n_911;
reg cadence_register_n_912;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_912 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_912 <= T_9_8_;
    end
 end
 assign n_912 = cadence_register_n_912;
reg cadence_register_n_913;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_913 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_913 <= sub_890_40_n_169;
    end
 end
 assign n_913 = cadence_register_n_913;
reg cadence_register_n_914;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_914 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_914 <= sub_890_40_n_184;
    end
 end
 assign n_914 = cadence_register_n_914;
reg cadence_register_n_915;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_915 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_915 <= sub_890_40_n_34;
    end
 end
 assign n_915 = cadence_register_n_915;
reg cadence_register_n_916;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_916 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_916 <= sub_890_40_n_33;
    end
 end
 assign n_916 = cadence_register_n_916;
reg cadence_register_n_917;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_917 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_917 <= R_10_21_;
    end
 end
 assign n_917 = cadence_register_n_917;
reg cadence_register_n_918;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_918 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_918 <= R_10_18_;
    end
 end
 assign n_918 = cadence_register_n_918;
reg cadence_register_n_919;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_919 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_919 <= sub_890_40_n_109;
    end
 end
 assign n_919 = cadence_register_n_919;
reg cadence_register_n_920;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_920 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_920 <= sub_890_40_n_26;
    end
 end
 assign n_920 = cadence_register_n_920;
reg cadence_register_n_921;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_921 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_921 <= R_10_14_;
    end
 end
 assign n_921 = cadence_register_n_921;
reg cadence_register_n_922;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_922 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_922 <= sub_890_40_n_100;
    end
 end
 assign n_922 = cadence_register_n_922;
reg cadence_register_n_923;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_923 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_923 <= R_10_19_;
    end
 end
 assign n_923 = cadence_register_n_923;
reg cadence_register_n_924;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_924 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_924 <= R_10_8_;
    end
 end
 assign n_924 = cadence_register_n_924;
reg cadence_register_n_925;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_925 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_925 <= sub_890_40_n_8;
    end
 end
 assign n_925 = cadence_register_n_925;
reg cadence_register_n_926;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_926 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_926 <= T_9_12_;
    end
 end
 assign n_926 = cadence_register_n_926;
reg cadence_register_n_927;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_927 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_927 <= sub_890_40_n_66;
    end
 end
 assign n_927 = cadence_register_n_927;
reg cadence_register_n_928;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_928 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_928 <= sub_890_40_n_126;
    end
 end
 assign n_928 = cadence_register_n_928;
reg cadence_register_n_929;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_929 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_929 <= T_9_9_;
    end
 end
 assign n_929 = cadence_register_n_929;
reg cadence_register_n_930;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_930 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_930 <= R_10_9_;
    end
 end
 assign n_930 = cadence_register_n_930;
reg cadence_register_n_931;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_931 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_931 <= T_9_10_;
    end
 end
 assign n_931 = cadence_register_n_931;
reg cadence_register_n_932;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_932 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_932 <= sub_890_40_n_19;
    end
 end
 assign n_932 = cadence_register_n_932;
reg cadence_register_n_933;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_933 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_933 <= T_9_6_;
    end
 end
 assign n_933 = cadence_register_n_933;
reg cadence_register_n_934;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_934 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_934 <= R_10_7_;
    end
 end
 assign n_934 = cadence_register_n_934;
reg cadence_register_n_935;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_935 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_935 <= T_9_5_;
    end
 end
 assign n_935 = cadence_register_n_935;
reg cadence_register_n_936;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_936 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_936 <= R_10_20_;
    end
 end
 assign n_936 = cadence_register_n_936;
reg cadence_register_n_937;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_937 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_937 <= sub_890_40_n_111;
    end
 end
 assign n_937 = cadence_register_n_937;
reg cadence_register_n_938;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_938 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_938 <= R_10_15_;
    end
 end
 assign n_938 = cadence_register_n_938;
reg cadence_register_n_939;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_939 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_939 <= sub_890_40_n_25;
    end
 end
 assign n_939 = cadence_register_n_939;
reg cadence_register_n_940;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_940 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_940 <= R_10_11_;
    end
 end
 assign n_940 = cadence_register_n_940;
reg cadence_register_n_941;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_941 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_941 <= sub_890_40_n_22;
    end
 end
 assign n_941 = cadence_register_n_941;
reg cadence_register_n_942;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_942 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_942 <= n_589;
    end
 end
 assign n_942 = cadence_register_n_942;
reg cadence_register_n_943;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_943 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_943 <= R_10_6_;
    end
 end
 assign n_943 = cadence_register_n_943;
reg cadence_register_n_944;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_944 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_944 <= R_10_12_;
    end
 end
 assign n_944 = cadence_register_n_944;
reg cadence_register_n_945;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_945 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_945 <= R_10_16_;
    end
 end
 assign n_945 = cadence_register_n_945;
reg cadence_register_n_946;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_946 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_946 <= sub_890_40_n_27;
    end
 end
 assign n_946 = cadence_register_n_946;
reg cadence_register_n_947;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_947 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_947 <= sub_890_40_n_119;
    end
 end
 assign n_947 = cadence_register_n_947;
reg cadence_register_n_948;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_948 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_948 <= R_10_0_;
    end
 end
 assign n_948 = cadence_register_n_948;
reg cadence_register_n_949;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_949 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_949 <= T_9_2_;
    end
 end
 assign n_949 = cadence_register_n_949;
reg cadence_register_n_950;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_950 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_950 <= n_592;
    end
 end
 assign n_950 = cadence_register_n_950;
reg cadence_register_n_951;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_951 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_951 <= n_590;
    end
 end
 assign n_951 = cadence_register_n_951;
reg cadence_register_n_952;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_952 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_952 <= T_9_4_;
    end
 end
 assign n_952 = cadence_register_n_952;
reg cadence_register_n_953;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_953 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_953 <= R_10_2_;
    end
 end
 assign n_953 = cadence_register_n_953;
reg cadence_register_n_954;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_954 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_954 <= R_10_3_;
    end
 end
 assign n_954 = cadence_register_n_954;
reg cadence_register_n_955;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_955 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_955 <= R_10_13_;
    end
 end
 assign n_955 = cadence_register_n_955;
reg cadence_register_n_956;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_956 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_956 <= sub_890_40_n_5;
    end
 end
 assign n_956 = cadence_register_n_956;
reg cadence_register_n_957;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_957 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_957 <= sub_890_40_n_120;
    end
 end
 assign n_957 = cadence_register_n_957;
reg cadence_register_n_958;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_958 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_958 <= sub_890_40_n_73;
    end
 end
 assign n_958 = cadence_register_n_958;
reg cadence_register_n_959;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_959 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_959 <= sub_890_40_n_83;
    end
 end
 assign n_959 = cadence_register_n_959;
reg cadence_register_n_960;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_960 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_960 <= R_10_5_;
    end
 end
 assign n_960 = cadence_register_n_960;
reg cadence_register_n_961;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_961 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_961 <= sub_890_40_n_182;
    end
 end
 assign n_961 = cadence_register_n_961;
reg cadence_register_n_962;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_962 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_962 <= sub_890_40_n_180;
    end
 end
 assign n_962 = cadence_register_n_962;
reg cadence_register_n_963;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_963 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_963 <= sub_890_40_n_116;
    end
 end
 assign n_963 = cadence_register_n_963;
reg cadence_register_n_964;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_964 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_964 <= n_593;
    end
 end
 assign n_964 = cadence_register_n_964;
reg cadence_register_n_965;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_965 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_965 <= n_198;
    end
 end
 assign n_965 = cadence_register_n_965;
reg cadence_register_n_966;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_966 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_966 <= R_14_1_;
    end
 end
 assign n_966 = cadence_register_n_966;
reg cadence_register_n_967;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_967 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_967 <= R_14_3_;
    end
 end
 assign n_967 = cadence_register_n_967;
reg cadence_register_n_968;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_968 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_968 <= R_14_8_;
    end
 end
 assign n_968 = cadence_register_n_968;
reg cadence_register_n_969;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_969 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_969 <= R_14_2_;
    end
 end
 assign n_969 = cadence_register_n_969;
reg cadence_register_n_970;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_970 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_970 <= R_14_9_;
    end
 end
 assign n_970 = cadence_register_n_970;
reg cadence_register_n_971;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_971 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_971 <= R_14_5_;
    end
 end
 assign n_971 = cadence_register_n_971;
reg cadence_register_n_972;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_972 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_972 <= R_14_13_;
    end
 end
 assign n_972 = cadence_register_n_972;
reg cadence_register_n_973;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_973 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_973 <= R_14_12_;
    end
 end
 assign n_973 = cadence_register_n_973;
reg cadence_register_n_974;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_974 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_974 <= T_14_11_;
    end
 end
 assign n_974 = cadence_register_n_974;
reg cadence_register_n_975;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_975 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_975 <= T_14_17_;
    end
 end
 assign n_975 = cadence_register_n_975;
reg cadence_register_n_976;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_976 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_976 <= T_14_32_;
    end
 end
 assign n_976 = cadence_register_n_976;
reg cadence_register_n_977;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_977 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_977 <= R_14_6_;
    end
 end
 assign n_977 = cadence_register_n_977;
reg cadence_register_n_978;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_978 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_978 <= R_14_7_;
    end
 end
 assign n_978 = cadence_register_n_978;
reg cadence_register_n_979;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_979 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_979 <= R_14_0_;
    end
 end
 assign n_979 = cadence_register_n_979;
reg cadence_register_n_980;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_980 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_980 <= R_14_16_;
    end
 end
 assign n_980 = cadence_register_n_980;
reg cadence_register_n_981;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_981 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_981 <= n_197;
    end
 end
 assign n_981 = cadence_register_n_981;
reg cadence_register_n_982;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_982 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_982 <= n_208;
    end
 end
 assign n_982 = cadence_register_n_982;
reg cadence_register_n_983;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_983 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_983 <= T_14_15_;
    end
 end
 assign n_983 = cadence_register_n_983;
reg cadence_register_n_984;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_984 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_984 <= R_14_10_;
    end
 end
 assign n_984 = cadence_register_n_984;
reg cadence_register_n_985;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_985 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_985 <= R_14_4_;
    end
 end
 assign n_985 = cadence_register_n_985;
reg cadence_register_n_986;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_986 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_986 <= R_14_14_;
    end
 end
 assign n_986 = cadence_register_n_986;
reg cadence_register_n_987;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_987 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_987 <= R_19_4_;
    end
 end
 assign n_987 = cadence_register_n_987;
reg cadence_register_n_988;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_988 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_988 <= sub_620_51_n_9;
    end
 end
 assign n_988 = cadence_register_n_988;
reg cadence_register_n_989;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_989 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_989 <= R_19_5_;
    end
 end
 assign n_989 = cadence_register_n_989;
reg cadence_register_n_990;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_990 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_990 <= sub_620_51_n_1;
    end
 end
 assign n_990 = cadence_register_n_990;
reg cadence_register_n_991;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_991 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_991 <= sub_620_51_n_28;
    end
 end
 assign n_991 = cadence_register_n_991;
reg cadence_register_n_992;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_992 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_992 <= R_19_11_;
    end
 end
 assign n_992 = cadence_register_n_992;
reg cadence_register_n_993;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_993 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_993 <= sub_620_51_n_52;
    end
 end
 assign n_993 = cadence_register_n_993;
reg cadence_register_n_994;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_994 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_994 <= R_19_10_;
    end
 end
 assign n_994 = cadence_register_n_994;
reg cadence_register_n_995;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_995 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_995 <= R_19_12_;
    end
 end
 assign n_995 = cadence_register_n_995;
reg cadence_register_n_996;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_996 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_996 <= R_19_8_;
    end
 end
 assign n_996 = cadence_register_n_996;
reg cadence_register_n_997;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_997 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_997 <= sub_620_51_n_42;
    end
 end
 assign n_997 = cadence_register_n_997;
reg cadence_register_n_998;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_998 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_998 <= sub_620_51_n_44;
    end
 end
 assign n_998 = cadence_register_n_998;
reg cadence_register_n_999;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_999 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_999 <= R_19_7_;
    end
 end
 assign n_999 = cadence_register_n_999;
reg cadence_register_n_1000;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1000 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1000 <= R_19_1_;
    end
 end
 assign n_1000 = cadence_register_n_1000;
reg cadence_register_n_1001;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1001 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1001 <= sub_620_51_n_46;
    end
 end
 assign n_1001 = cadence_register_n_1001;
reg cadence_register_n_1002;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1002 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1002 <= sub_620_51_n_5;
    end
 end
 assign n_1002 = cadence_register_n_1002;
reg cadence_register_n_1003;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1003 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1003 <= R_19_2_;
    end
 end
 assign n_1003 = cadence_register_n_1003;
reg cadence_register_n_1004;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1004 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1004 <= R_19_3_;
    end
 end
 assign n_1004 = cadence_register_n_1004;
reg cadence_register_n_1005;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1005 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1005 <= sub_620_51_n_27;
    end
 end
 assign n_1005 = cadence_register_n_1005;
reg cadence_register_n_1006;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1006 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1006 <= sub_620_51_n_53;
    end
 end
 assign n_1006 = cadence_register_n_1006;
reg cadence_register_n_1007;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1007 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1007 <= sub_620_51_n_37;
    end
 end
 assign n_1007 = cadence_register_n_1007;
reg cadence_register_n_1008;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1008 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1008 <= R_19_0_;
    end
 end
 assign n_1008 = cadence_register_n_1008;
reg cadence_register_n_1009;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1009 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1009 <= sub_620_51_n_8;
    end
 end
 assign n_1009 = cadence_register_n_1009;
reg cadence_register_n_1010;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1010 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1010 <= sub_620_51_n_40;
    end
 end
 assign n_1010 = cadence_register_n_1010;
reg cadence_register_n_1011;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1011 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1011 <= sub_620_51_n_30;
    end
 end
 assign n_1011 = cadence_register_n_1011;
reg cadence_register_n_1012;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1012 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1012 <= sub_620_51_n_6;
    end
 end
 assign n_1012 = cadence_register_n_1012;
reg cadence_register_n_1013;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1013 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1013 <= R_19_6_;
    end
 end
 assign n_1013 = cadence_register_n_1013;
reg cadence_register_n_1014;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1014 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1014 <= sub_620_51_n_25;
    end
 end
 assign n_1014 = cadence_register_n_1014;
reg cadence_register_n_1015;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1015 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1015 <= sub_620_51_n_7;
    end
 end
 assign n_1015 = cadence_register_n_1015;
reg cadence_register_n_1016;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1016 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1016 <= R_19_9_;
    end
 end
 assign n_1016 = cadence_register_n_1016;
reg cadence_register_n_1017;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1017 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1017 <= in2[23];
    end
 end
 assign n_1017 = cadence_register_n_1017;
reg cadence_register_n_1018;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1018 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1018 <= in2[21];
    end
 end
 assign n_1018 = cadence_register_n_1018;
reg cadence_register_n_1019;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1019 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1019 <= sub_470_56_n_17;
    end
 end
 assign n_1019 = cadence_register_n_1019;
reg cadence_register_n_1020;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1020 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1020 <= T_24_2_;
    end
 end
 assign n_1020 = cadence_register_n_1020;
reg cadence_register_n_1021;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1021 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1021 <= T_24_32_;
    end
 end
 assign n_1021 = cadence_register_n_1021;
reg cadence_register_n_1022;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1022 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1022 <= n_42;
    end
 end
 assign n_1022 = cadence_register_n_1022;
reg cadence_register_n_1023;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1023 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1023 <= n_36;
    end
 end
 assign n_1023 = cadence_register_n_1023;
reg cadence_register_n_1024;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1024 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1024 <= in2[19];
    end
 end
 assign n_1024 = cadence_register_n_1024;
reg cadence_register_n_1025;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1025 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1025 <= in1[12];
    end
 end
 assign n_1025 = cadence_register_n_1025;
reg cadence_register_n_1026;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1026 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1026 <= n_1025;
    end
 end
 assign n_1026 = cadence_register_n_1026;
reg cadence_register_n_1027;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1027 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1027 <= n_1026;
    end
 end
 assign n_1027 = cadence_register_n_1027;
reg cadence_register_n_1028;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1028 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1028 <= n_1027;
    end
 end
 assign n_1028 = cadence_register_n_1028;
reg cadence_register_n_1029;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1029 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1029 <= n_1028;
    end
 end
 assign n_1029 = cadence_register_n_1029;
reg cadence_register_n_1030;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1030 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1030 <= in1[18];
    end
 end
 assign n_1030 = cadence_register_n_1030;
reg cadence_register_n_1031;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1031 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1031 <= n_1030;
    end
 end
 assign n_1031 = cadence_register_n_1031;
reg cadence_register_n_1032;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1032 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1032 <= n_1031;
    end
 end
 assign n_1032 = cadence_register_n_1032;
reg cadence_register_n_1033;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1033 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1033 <= n_1032;
    end
 end
 assign n_1033 = cadence_register_n_1033;
reg cadence_register_n_1034;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1034 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1034 <= n_1033;
    end
 end
 assign n_1034 = cadence_register_n_1034;
reg cadence_register_n_1035;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1035 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1035 <= in2[5];
    end
 end
 assign n_1035 = cadence_register_n_1035;
reg cadence_register_n_1036;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1036 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1036 <= n_1035;
    end
 end
 assign n_1036 = cadence_register_n_1036;
reg cadence_register_n_1037;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1037 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1037 <= n_1036;
    end
 end
 assign n_1037 = cadence_register_n_1037;
reg cadence_register_n_1038;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1038 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1038 <= n_1037;
    end
 end
 assign n_1038 = cadence_register_n_1038;
reg cadence_register_n_1039;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1039 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1039 <= sub_1010_35_n_83;
    end
 end
 assign n_1039 = cadence_register_n_1039;
reg cadence_register_n_1040;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1040 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1040 <= n_1039;
    end
 end
 assign n_1040 = cadence_register_n_1040;
reg cadence_register_n_1041;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1041 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1041 <= n_1040;
    end
 end
 assign n_1041 = cadence_register_n_1041;
reg cadence_register_n_1042;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1042 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1042 <= n_1041;
    end
 end
 assign n_1042 = cadence_register_n_1042;
reg cadence_register_n_1043;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1043 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1043 <= n_35;
    end
 end
 assign n_1043 = cadence_register_n_1043;
reg cadence_register_n_1044;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1044 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1044 <= n_529;
    end
 end
 assign n_1044 = cadence_register_n_1044;
reg cadence_register_n_1045;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1045 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1045 <= n_1044;
    end
 end
 assign n_1045 = cadence_register_n_1045;
reg cadence_register_n_1046;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1046 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1046 <= n_1045;
    end
 end
 assign n_1046 = cadence_register_n_1046;
reg cadence_register_n_1047;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1047 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1047 <= n_1046;
    end
 end
 assign n_1047 = cadence_register_n_1047;
reg cadence_register_n_1048;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1048 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1048 <= in1[5];
    end
 end
 assign n_1048 = cadence_register_n_1048;
reg cadence_register_n_1049;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1049 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1049 <= n_1048;
    end
 end
 assign n_1049 = cadence_register_n_1049;
reg cadence_register_n_1050;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1050 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1050 <= n_1049;
    end
 end
 assign n_1050 = cadence_register_n_1050;
reg cadence_register_n_1051;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1051 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1051 <= n_1050;
    end
 end
 assign n_1051 = cadence_register_n_1051;
reg cadence_register_n_1052;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1052 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1052 <= n_1051;
    end
 end
 assign n_1052 = cadence_register_n_1052;
reg cadence_register_n_1053;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1053 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1053 <= n_30;
    end
 end
 assign n_1053 = cadence_register_n_1053;
reg cadence_register_n_1054;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1054 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1054 <= T_24_6_;
    end
 end
 assign n_1054 = cadence_register_n_1054;
reg cadence_register_n_1055;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1055 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1055 <= in2[17];
    end
 end
 assign n_1055 = cadence_register_n_1055;
reg cadence_register_n_1056;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1056 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1056 <= n_1055;
    end
 end
 assign n_1056 = cadence_register_n_1056;
reg cadence_register_n_1057;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1057 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1057 <= in2[22];
    end
 end
 assign n_1057 = cadence_register_n_1057;
reg cadence_register_n_1058;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1058 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1058 <= in1[24];
    end
 end
 assign n_1058 = cadence_register_n_1058;
reg cadence_register_n_1059;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1059 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1059 <= n_1058;
    end
 end
 assign n_1059 = cadence_register_n_1059;
reg cadence_register_n_1060;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1060 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1060 <= n_1059;
    end
 end
 assign n_1060 = cadence_register_n_1060;
reg cadence_register_n_1061;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1061 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1061 <= n_1060;
    end
 end
 assign n_1061 = cadence_register_n_1061;
reg cadence_register_n_1062;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1062 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1062 <= n_1061;
    end
 end
 assign n_1062 = cadence_register_n_1062;
reg cadence_register_n_1063;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1063 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1063 <= sub_1040_34_n_62;
    end
 end
 assign n_1063 = cadence_register_n_1063;
reg cadence_register_n_1064;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1064 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1064 <= in1[11];
    end
 end
 assign n_1064 = cadence_register_n_1064;
reg cadence_register_n_1065;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1065 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1065 <= n_1064;
    end
 end
 assign n_1065 = cadence_register_n_1065;
reg cadence_register_n_1066;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1066 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1066 <= n_1065;
    end
 end
 assign n_1066 = cadence_register_n_1066;
reg cadence_register_n_1067;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1067 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1067 <= n_1066;
    end
 end
 assign n_1067 = cadence_register_n_1067;
reg cadence_register_n_1068;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1068 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1068 <= n_1067;
    end
 end
 assign n_1068 = cadence_register_n_1068;
reg cadence_register_n_1069;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1069 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1069 <= in2[11];
    end
 end
 assign n_1069 = cadence_register_n_1069;
reg cadence_register_n_1070;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1070 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1070 <= n_1069;
    end
 end
 assign n_1070 = cadence_register_n_1070;
reg cadence_register_n_1071;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1071 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1071 <= n_1070;
    end
 end
 assign n_1071 = cadence_register_n_1071;
reg cadence_register_n_1072;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1072 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1072 <= sub_830_44_n_72;
    end
 end
 assign n_1072 = cadence_register_n_1072;
reg cadence_register_n_1073;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1073 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1073 <= n_1072;
    end
 end
 assign n_1073 = cadence_register_n_1073;
reg cadence_register_n_1074;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1074 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1074 <= n_1073;
    end
 end
 assign n_1074 = cadence_register_n_1074;
reg cadence_register_n_1075;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1075 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1075 <= T_11_0_;
    end
 end
 assign n_1075 = cadence_register_n_1075;
reg cadence_register_n_1076;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1076 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1076 <= n_1075;
    end
 end
 assign n_1076 = cadence_register_n_1076;
reg cadence_register_n_1077;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1077 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1077 <= n_1076;
    end
 end
 assign n_1077 = cadence_register_n_1077;
reg cadence_register_n_1078;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1078 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1078 <= n_31;
    end
 end
 assign n_1078 = cadence_register_n_1078;
reg cadence_register_n_1079;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1079 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1079 <= n_38;
    end
 end
 assign n_1079 = cadence_register_n_1079;
reg cadence_register_n_1080;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1080 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1080 <= T_24_7_;
    end
 end
 assign n_1080 = cadence_register_n_1080;
reg cadence_register_n_1081;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1081 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1081 <= T_24_1_;
    end
 end
 assign n_1081 = cadence_register_n_1081;
reg cadence_register_n_1082;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1082 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1082 <= n_33;
    end
 end
 assign n_1082 = cadence_register_n_1082;
reg cadence_register_n_1083;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1083 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1083 <= in2[16];
    end
 end
 assign n_1083 = cadence_register_n_1083;
reg cadence_register_n_1084;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1084 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1084 <= n_1083;
    end
 end
 assign n_1084 = cadence_register_n_1084;
reg cadence_register_n_1085;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1085 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1085 <= in1[26];
    end
 end
 assign n_1085 = cadence_register_n_1085;
reg cadence_register_n_1086;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1086 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1086 <= n_1085;
    end
 end
 assign n_1086 = cadence_register_n_1086;
reg cadence_register_n_1087;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1087 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1087 <= n_1086;
    end
 end
 assign n_1087 = cadence_register_n_1087;
reg cadence_register_n_1088;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1088 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1088 <= n_1087;
    end
 end
 assign n_1088 = cadence_register_n_1088;
reg cadence_register_n_1089;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1089 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1089 <= n_1088;
    end
 end
 assign n_1089 = cadence_register_n_1089;
reg cadence_register_n_1090;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1090 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1090 <= in1[15];
    end
 end
 assign n_1090 = cadence_register_n_1090;
reg cadence_register_n_1091;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1091 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1091 <= n_1090;
    end
 end
 assign n_1091 = cadence_register_n_1091;
reg cadence_register_n_1092;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1092 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1092 <= n_1091;
    end
 end
 assign n_1092 = cadence_register_n_1092;
reg cadence_register_n_1093;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1093 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1093 <= n_1092;
    end
 end
 assign n_1093 = cadence_register_n_1093;
reg cadence_register_n_1094;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1094 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1094 <= n_1093;
    end
 end
 assign n_1094 = cadence_register_n_1094;
reg cadence_register_n_1095;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1095 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1095 <= in1[6];
    end
 end
 assign n_1095 = cadence_register_n_1095;
reg cadence_register_n_1096;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1096 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1096 <= n_1095;
    end
 end
 assign n_1096 = cadence_register_n_1096;
reg cadence_register_n_1097;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1097 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1097 <= n_1096;
    end
 end
 assign n_1097 = cadence_register_n_1097;
reg cadence_register_n_1098;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1098 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1098 <= n_1097;
    end
 end
 assign n_1098 = cadence_register_n_1098;
reg cadence_register_n_1099;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1099 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1099 <= n_1098;
    end
 end
 assign n_1099 = cadence_register_n_1099;
reg cadence_register_n_1100;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1100 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1100 <= in1[2];
    end
 end
 assign n_1100 = cadence_register_n_1100;
reg cadence_register_n_1101;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1101 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1101 <= n_1100;
    end
 end
 assign n_1101 = cadence_register_n_1101;
reg cadence_register_n_1102;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1102 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1102 <= n_1101;
    end
 end
 assign n_1102 = cadence_register_n_1102;
reg cadence_register_n_1103;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1103 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1103 <= n_1102;
    end
 end
 assign n_1103 = cadence_register_n_1103;
reg cadence_register_n_1104;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1104 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1104 <= n_1103;
    end
 end
 assign n_1104 = cadence_register_n_1104;
reg cadence_register_n_1105;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1105 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1105 <= T_16_0_;
    end
 end
 assign n_1105 = cadence_register_n_1105;
reg cadence_register_n_1106;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1106 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1106 <= n_1105;
    end
 end
 assign n_1106 = cadence_register_n_1106;
reg cadence_register_n_1107;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1107 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1107 <= n_29;
    end
 end
 assign n_1107 = cadence_register_n_1107;
reg cadence_register_n_1108;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1108 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1108 <= n_34;
    end
 end
 assign n_1108 = cadence_register_n_1108;
reg cadence_register_n_1109;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1109 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1109 <= in2[20];
    end
 end
 assign n_1109 = cadence_register_n_1109;
reg cadence_register_n_1110;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1110 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1110 <= in2[15];
    end
 end
 assign n_1110 = cadence_register_n_1110;
reg cadence_register_n_1111;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1111 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1111 <= n_1110;
    end
 end
 assign n_1111 = cadence_register_n_1111;
reg cadence_register_n_1112;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1112 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1112 <= in1[3];
    end
 end
 assign n_1112 = cadence_register_n_1112;
reg cadence_register_n_1113;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1113 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1113 <= n_1112;
    end
 end
 assign n_1113 = cadence_register_n_1113;
reg cadence_register_n_1114;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1114 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1114 <= n_1113;
    end
 end
 assign n_1114 = cadence_register_n_1114;
reg cadence_register_n_1115;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1115 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1115 <= n_1114;
    end
 end
 assign n_1115 = cadence_register_n_1115;
reg cadence_register_n_1116;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1116 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1116 <= n_1115;
    end
 end
 assign n_1116 = cadence_register_n_1116;
reg cadence_register_n_1117;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1117 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1117 <= n_37;
    end
 end
 assign n_1117 = cadence_register_n_1117;
reg cadence_register_n_1118;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1118 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1118 <= T_15_0_;
    end
 end
 assign n_1118 = cadence_register_n_1118;
reg cadence_register_n_1119;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1119 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1119 <= n_1118;
    end
 end
 assign n_1119 = cadence_register_n_1119;
reg cadence_register_n_1120;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1120 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1120 <= in2[18];
    end
 end
 assign n_1120 = cadence_register_n_1120;
reg cadence_register_n_1121;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1121 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1121 <= n_1120;
    end
 end
 assign n_1121 = cadence_register_n_1121;
reg cadence_register_n_1122;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1122 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1122 <= in2[4];
    end
 end
 assign n_1122 = cadence_register_n_1122;
reg cadence_register_n_1123;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1123 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1123 <= n_1122;
    end
 end
 assign n_1123 = cadence_register_n_1123;
reg cadence_register_n_1124;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1124 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1124 <= n_1123;
    end
 end
 assign n_1124 = cadence_register_n_1124;
reg cadence_register_n_1125;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1125 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1125 <= n_1124;
    end
 end
 assign n_1125 = cadence_register_n_1125;
reg cadence_register_n_1126;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1126 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1126 <= n_1125;
    end
 end
 assign n_1126 = cadence_register_n_1126;
reg cadence_register_n_1127;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1127 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1127 <= sub_620_51_n_36;
    end
 end
 assign n_1127 = cadence_register_n_1127;
reg cadence_register_n_1128;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1128 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1128 <= n_1127;
    end
 end
 assign n_1128 = cadence_register_n_1128;
reg cadence_register_n_1129;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1129 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1129 <= sub_1040_34_n_93;
    end
 end
 assign n_1129 = cadence_register_n_1129;
reg cadence_register_n_1130;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1130 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1130 <= n_1129;
    end
 end
 assign n_1130 = cadence_register_n_1130;
reg cadence_register_n_1131;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1131 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1131 <= n_1130;
    end
 end
 assign n_1131 = cadence_register_n_1131;
reg cadence_register_n_1132;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1132 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1132 <= n_1131;
    end
 end
 assign n_1132 = cadence_register_n_1132;
reg cadence_register_n_1133;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1133 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1133 <= T_18_0_;
    end
 end
 assign n_1133 = cadence_register_n_1133;
reg cadence_register_n_1134;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1134 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1134 <= n_1133;
    end
 end
 assign n_1134 = cadence_register_n_1134;
reg cadence_register_n_1135;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1135 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1135 <= in1[16];
    end
 end
 assign n_1135 = cadence_register_n_1135;
reg cadence_register_n_1136;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1136 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1136 <= n_1135;
    end
 end
 assign n_1136 = cadence_register_n_1136;
reg cadence_register_n_1137;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1137 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1137 <= n_1136;
    end
 end
 assign n_1137 = cadence_register_n_1137;
reg cadence_register_n_1138;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1138 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1138 <= n_1137;
    end
 end
 assign n_1138 = cadence_register_n_1138;
reg cadence_register_n_1139;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1139 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1139 <= n_1138;
    end
 end
 assign n_1139 = cadence_register_n_1139;
reg cadence_register_n_1140;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1140 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1140 <= in2[7];
    end
 end
 assign n_1140 = cadence_register_n_1140;
reg cadence_register_n_1141;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1141 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1141 <= n_1140;
    end
 end
 assign n_1141 = cadence_register_n_1141;
reg cadence_register_n_1142;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1142 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1142 <= n_1141;
    end
 end
 assign n_1142 = cadence_register_n_1142;
reg cadence_register_n_1143;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1143 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1143 <= n_1142;
    end
 end
 assign n_1143 = cadence_register_n_1143;
reg cadence_register_n_1144;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1144 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1144 <= in2[13];
    end
 end
 assign n_1144 = cadence_register_n_1144;
reg cadence_register_n_1145;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1145 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1145 <= n_1144;
    end
 end
 assign n_1145 = cadence_register_n_1145;
reg cadence_register_n_1146;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1146 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1146 <= n_1145;
    end
 end
 assign n_1146 = cadence_register_n_1146;
reg cadence_register_n_1147;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1147 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1147 <= sub_950_37_n_68;
    end
 end
 assign n_1147 = cadence_register_n_1147;
reg cadence_register_n_1148;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1148 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1148 <= n_1147;
    end
 end
 assign n_1148 = cadence_register_n_1148;
reg cadence_register_n_1149;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1149 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1149 <= n_1148;
    end
 end
 assign n_1149 = cadence_register_n_1149;
reg cadence_register_n_1150;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1150 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1150 <= n_1149;
    end
 end
 assign n_1150 = cadence_register_n_1150;
reg cadence_register_n_1151;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1151 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1151 <= sub_770_46_n_56;
    end
 end
 assign n_1151 = cadence_register_n_1151;
reg cadence_register_n_1152;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1152 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1152 <= n_1151;
    end
 end
 assign n_1152 = cadence_register_n_1152;
reg cadence_register_n_1153;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1153 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1153 <= n_1152;
    end
 end
 assign n_1153 = cadence_register_n_1153;
reg cadence_register_n_1154;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1154 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1154 <= T_13_0_;
    end
 end
 assign n_1154 = cadence_register_n_1154;
reg cadence_register_n_1155;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1155 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1155 <= n_1154;
    end
 end
 assign n_1155 = cadence_register_n_1155;
reg cadence_register_n_1156;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1156 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1156 <= n_1155;
    end
 end
 assign n_1156 = cadence_register_n_1156;
reg cadence_register_n_1157;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1157 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1157 <= T_7_0_;
    end
 end
 assign n_1157 = cadence_register_n_1157;
reg cadence_register_n_1158;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1158 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1158 <= n_1157;
    end
 end
 assign n_1158 = cadence_register_n_1158;
reg cadence_register_n_1159;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1159 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1159 <= n_1158;
    end
 end
 assign n_1159 = cadence_register_n_1159;
reg cadence_register_n_1160;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1160 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1160 <= n_1159;
    end
 end
 assign n_1160 = cadence_register_n_1160;
reg cadence_register_n_1161;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1161 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1161 <= in1[9];
    end
 end
 assign n_1161 = cadence_register_n_1161;
reg cadence_register_n_1162;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1162 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1162 <= n_1161;
    end
 end
 assign n_1162 = cadence_register_n_1162;
reg cadence_register_n_1163;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1163 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1163 <= n_1162;
    end
 end
 assign n_1163 = cadence_register_n_1163;
reg cadence_register_n_1164;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1164 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1164 <= n_1163;
    end
 end
 assign n_1164 = cadence_register_n_1164;
reg cadence_register_n_1165;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1165 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1165 <= n_1164;
    end
 end
 assign n_1165 = cadence_register_n_1165;
reg cadence_register_n_1166;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1166 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1166 <= in1[7];
    end
 end
 assign n_1166 = cadence_register_n_1166;
reg cadence_register_n_1167;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1167 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1167 <= n_1166;
    end
 end
 assign n_1167 = cadence_register_n_1167;
reg cadence_register_n_1168;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1168 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1168 <= n_1167;
    end
 end
 assign n_1168 = cadence_register_n_1168;
reg cadence_register_n_1169;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1169 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1169 <= n_1168;
    end
 end
 assign n_1169 = cadence_register_n_1169;
reg cadence_register_n_1170;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1170 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1170 <= n_1169;
    end
 end
 assign n_1170 = cadence_register_n_1170;
reg cadence_register_n_1171;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1171 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1171 <= in1[17];
    end
 end
 assign n_1171 = cadence_register_n_1171;
reg cadence_register_n_1172;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1172 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1172 <= n_1171;
    end
 end
 assign n_1172 = cadence_register_n_1172;
reg cadence_register_n_1173;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1173 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1173 <= n_1172;
    end
 end
 assign n_1173 = cadence_register_n_1173;
reg cadence_register_n_1174;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1174 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1174 <= n_1173;
    end
 end
 assign n_1174 = cadence_register_n_1174;
reg cadence_register_n_1175;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1175 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1175 <= n_1174;
    end
 end
 assign n_1175 = cadence_register_n_1175;
reg cadence_register_n_1176;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1176 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1176 <= in1[22];
    end
 end
 assign n_1176 = cadence_register_n_1176;
reg cadence_register_n_1177;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1177 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1177 <= n_1176;
    end
 end
 assign n_1177 = cadence_register_n_1177;
reg cadence_register_n_1178;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1178 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1178 <= n_1177;
    end
 end
 assign n_1178 = cadence_register_n_1178;
reg cadence_register_n_1179;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1179 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1179 <= n_1178;
    end
 end
 assign n_1179 = cadence_register_n_1179;
reg cadence_register_n_1180;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1180 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1180 <= n_1179;
    end
 end
 assign n_1180 = cadence_register_n_1180;
reg cadence_register_n_1181;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1181 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1181 <= in1[14];
    end
 end
 assign n_1181 = cadence_register_n_1181;
reg cadence_register_n_1182;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1182 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1182 <= n_1181;
    end
 end
 assign n_1182 = cadence_register_n_1182;
reg cadence_register_n_1183;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1183 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1183 <= n_1182;
    end
 end
 assign n_1183 = cadence_register_n_1183;
reg cadence_register_n_1184;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1184 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1184 <= n_1183;
    end
 end
 assign n_1184 = cadence_register_n_1184;
reg cadence_register_n_1185;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1185 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1185 <= n_1184;
    end
 end
 assign n_1185 = cadence_register_n_1185;
reg cadence_register_n_1186;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1186 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1186 <= in2[14];
    end
 end
 assign n_1186 = cadence_register_n_1186;
reg cadence_register_n_1187;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1187 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1187 <= n_1186;
    end
 end
 assign n_1187 = cadence_register_n_1187;
reg cadence_register_n_1188;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1188 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1188 <= sub_740_47_n_57;
    end
 end
 assign n_1188 = cadence_register_n_1188;
reg cadence_register_n_1189;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1189 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1189 <= n_1188;
    end
 end
 assign n_1189 = cadence_register_n_1189;
reg cadence_register_n_1190;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1190 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1190 <= T_14_0_;
    end
 end
 assign n_1190 = cadence_register_n_1190;
reg cadence_register_n_1191;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1191 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1191 <= n_1190;
    end
 end
 assign n_1191 = cadence_register_n_1191;
reg cadence_register_n_1192;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1192 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1192 <= in2[8];
    end
 end
 assign n_1192 = cadence_register_n_1192;
reg cadence_register_n_1193;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1193 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1193 <= n_1192;
    end
 end
 assign n_1193 = cadence_register_n_1193;
reg cadence_register_n_1194;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1194 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1194 <= n_1193;
    end
 end
 assign n_1194 = cadence_register_n_1194;
reg cadence_register_n_1195;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1195 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1195 <= n_1194;
    end
 end
 assign n_1195 = cadence_register_n_1195;
reg cadence_register_n_1196;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1196 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1196 <= sub_920_38_n_57;
    end
 end
 assign n_1196 = cadence_register_n_1196;
reg cadence_register_n_1197;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1197 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1197 <= n_1196;
    end
 end
 assign n_1197 = cadence_register_n_1197;
reg cadence_register_n_1198;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1198 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1198 <= n_1197;
    end
 end
 assign n_1198 = cadence_register_n_1198;
reg cadence_register_n_1199;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1199 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1199 <= n_1198;
    end
 end
 assign n_1199 = cadence_register_n_1199;
reg cadence_register_n_1200;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1200 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1200 <= T_8_0_;
    end
 end
 assign n_1200 = cadence_register_n_1200;
reg cadence_register_n_1201;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1201 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1201 <= n_1200;
    end
 end
 assign n_1201 = cadence_register_n_1201;
reg cadence_register_n_1202;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1202 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1202 <= n_1201;
    end
 end
 assign n_1202 = cadence_register_n_1202;
reg cadence_register_n_1203;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1203 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1203 <= n_1202;
    end
 end
 assign n_1203 = cadence_register_n_1203;
reg cadence_register_n_1204;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1204 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1204 <= in2[10];
    end
 end
 assign n_1204 = cadence_register_n_1204;
reg cadence_register_n_1205;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1205 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1205 <= n_1204;
    end
 end
 assign n_1205 = cadence_register_n_1205;
reg cadence_register_n_1206;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1206 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1206 <= n_1205;
    end
 end
 assign n_1206 = cadence_register_n_1206;
reg cadence_register_n_1207;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1207 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1207 <= T_24_0_;
    end
 end
 assign n_1207 = cadence_register_n_1207;
reg cadence_register_n_1208;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1208 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1208 <= sub_860_43_n_70;
    end
 end
 assign n_1208 = cadence_register_n_1208;
reg cadence_register_n_1209;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1209 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1209 <= n_1208;
    end
 end
 assign n_1209 = cadence_register_n_1209;
reg cadence_register_n_1210;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1210 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1210 <= n_1209;
    end
 end
 assign n_1210 = cadence_register_n_1210;
reg cadence_register_n_1211;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1211 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1211 <= in1[20];
    end
 end
 assign n_1211 = cadence_register_n_1211;
reg cadence_register_n_1212;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1212 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1212 <= n_1211;
    end
 end
 assign n_1212 = cadence_register_n_1212;
reg cadence_register_n_1213;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1213 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1213 <= n_1212;
    end
 end
 assign n_1213 = cadence_register_n_1213;
reg cadence_register_n_1214;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1214 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1214 <= n_1213;
    end
 end
 assign n_1214 = cadence_register_n_1214;
reg cadence_register_n_1215;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1215 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1215 <= n_1214;
    end
 end
 assign n_1215 = cadence_register_n_1215;
reg cadence_register_n_1216;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1216 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1216 <= in1[8];
    end
 end
 assign n_1216 = cadence_register_n_1216;
reg cadence_register_n_1217;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1217 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1217 <= n_1216;
    end
 end
 assign n_1217 = cadence_register_n_1217;
reg cadence_register_n_1218;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1218 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1218 <= n_1217;
    end
 end
 assign n_1218 = cadence_register_n_1218;
reg cadence_register_n_1219;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1219 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1219 <= n_1218;
    end
 end
 assign n_1219 = cadence_register_n_1219;
reg cadence_register_n_1220;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1220 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1220 <= n_1219;
    end
 end
 assign n_1220 = cadence_register_n_1220;
reg cadence_register_n_1221;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1221 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1221 <= in2[6];
    end
 end
 assign n_1221 = cadence_register_n_1221;
reg cadence_register_n_1222;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1222 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1222 <= n_1221;
    end
 end
 assign n_1222 = cadence_register_n_1222;
reg cadence_register_n_1223;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1223 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1223 <= n_1222;
    end
 end
 assign n_1223 = cadence_register_n_1223;
reg cadence_register_n_1224;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1224 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1224 <= n_1223;
    end
 end
 assign n_1224 = cadence_register_n_1224;
reg cadence_register_n_1225;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1225 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1225 <= sub_980_36_n_68;
    end
 end
 assign n_1225 = cadence_register_n_1225;
reg cadence_register_n_1226;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1226 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1226 <= n_1225;
    end
 end
 assign n_1226 = cadence_register_n_1226;
reg cadence_register_n_1227;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1227 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1227 <= n_1226;
    end
 end
 assign n_1227 = cadence_register_n_1227;
reg cadence_register_n_1228;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1228 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1228 <= n_1227;
    end
 end
 assign n_1228 = cadence_register_n_1228;
reg cadence_register_n_1229;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1229 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1229 <= T_6_0_;
    end
 end
 assign n_1229 = cadence_register_n_1229;
reg cadence_register_n_1230;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1230 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1230 <= n_1229;
    end
 end
 assign n_1230 = cadence_register_n_1230;
reg cadence_register_n_1231;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1231 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1231 <= n_1230;
    end
 end
 assign n_1231 = cadence_register_n_1231;
reg cadence_register_n_1232;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1232 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1232 <= n_1231;
    end
 end
 assign n_1232 = cadence_register_n_1232;
reg cadence_register_n_1233;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1233 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1233 <= n_39;
    end
 end
 assign n_1233 = cadence_register_n_1233;
reg cadence_register_n_1234;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1234 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1234 <= in2[9];
    end
 end
 assign n_1234 = cadence_register_n_1234;
reg cadence_register_n_1235;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1235 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1235 <= n_1234;
    end
 end
 assign n_1235 = cadence_register_n_1235;
reg cadence_register_n_1236;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1236 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1236 <= n_1235;
    end
 end
 assign n_1236 = cadence_register_n_1236;
reg cadence_register_n_1237;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1237 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1237 <= n_1236;
    end
 end
 assign n_1237 = cadence_register_n_1237;
reg cadence_register_n_1238;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1238 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1238 <= sub_890_40_n_70;
    end
 end
 assign n_1238 = cadence_register_n_1238;
reg cadence_register_n_1239;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1239 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1239 <= n_1238;
    end
 end
 assign n_1239 = cadence_register_n_1239;
reg cadence_register_n_1240;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1240 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1240 <= n_1239;
    end
 end
 assign n_1240 = cadence_register_n_1240;
reg cadence_register_n_1241;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1241 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1241 <= in1[27];
    end
 end
 assign n_1241 = cadence_register_n_1241;
reg cadence_register_n_1242;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1242 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1242 <= n_1241;
    end
 end
 assign n_1242 = cadence_register_n_1242;
reg cadence_register_n_1243;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1243 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1243 <= n_1242;
    end
 end
 assign n_1243 = cadence_register_n_1243;
reg cadence_register_n_1244;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1244 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1244 <= n_1243;
    end
 end
 assign n_1244 = cadence_register_n_1244;
reg cadence_register_n_1245;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1245 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1245 <= n_1244;
    end
 end
 assign n_1245 = cadence_register_n_1245;
reg cadence_register_n_1246;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1246 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1246 <= in2[2];
    end
 end
 assign n_1246 = cadence_register_n_1246;
reg cadence_register_n_1247;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1247 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1247 <= n_1246;
    end
 end
 assign n_1247 = cadence_register_n_1247;
reg cadence_register_n_1248;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1248 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1248 <= n_1247;
    end
 end
 assign n_1248 = cadence_register_n_1248;
reg cadence_register_n_1249;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1249 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1249 <= n_1248;
    end
 end
 assign n_1249 = cadence_register_n_1249;
reg cadence_register_n_1250;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1250 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1250 <= n_1249;
    end
 end
 assign n_1250 = cadence_register_n_1250;
reg cadence_register_n_1251;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1251 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1251 <= sub_1100_32_n_96;
    end
 end
 assign n_1251 = cadence_register_n_1251;
reg cadence_register_n_1252;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1252 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1252 <= n_1251;
    end
 end
 assign n_1252 = cadence_register_n_1252;
reg cadence_register_n_1253;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1253 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1253 <= n_1252;
    end
 end
 assign n_1253 = cadence_register_n_1253;
reg cadence_register_n_1254;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1254 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1254 <= n_1253;
    end
 end
 assign n_1254 = cadence_register_n_1254;
reg cadence_register_n_1255;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1255 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1255 <= n_1254;
    end
 end
 assign n_1255 = cadence_register_n_1255;
reg cadence_register_n_1256;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1256 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1256 <= sub_680_49_n_51;
    end
 end
 assign n_1256 = cadence_register_n_1256;
reg cadence_register_n_1257;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1257 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1257 <= n_1256;
    end
 end
 assign n_1257 = cadence_register_n_1257;
reg cadence_register_n_1258;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1258 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1258 <= in1[13];
    end
 end
 assign n_1258 = cadence_register_n_1258;
reg cadence_register_n_1259;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1259 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1259 <= n_1258;
    end
 end
 assign n_1259 = cadence_register_n_1259;
reg cadence_register_n_1260;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1260 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1260 <= n_1259;
    end
 end
 assign n_1260 = cadence_register_n_1260;
reg cadence_register_n_1261;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1261 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1261 <= n_1260;
    end
 end
 assign n_1261 = cadence_register_n_1261;
reg cadence_register_n_1262;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1262 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1262 <= n_1261;
    end
 end
 assign n_1262 = cadence_register_n_1262;
reg cadence_register_n_1263;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1263 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1263 <= in2[12];
    end
 end
 assign n_1263 = cadence_register_n_1263;
reg cadence_register_n_1264;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1264 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1264 <= n_1263;
    end
 end
 assign n_1264 = cadence_register_n_1264;
reg cadence_register_n_1265;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1265 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1265 <= n_1264;
    end
 end
 assign n_1265 = cadence_register_n_1265;
reg cadence_register_n_1266;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1266 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1266 <= sub_800_45_n_58;
    end
 end
 assign n_1266 = cadence_register_n_1266;
reg cadence_register_n_1267;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1267 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1267 <= n_1266;
    end
 end
 assign n_1267 = cadence_register_n_1267;
reg cadence_register_n_1268;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1268 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1268 <= n_1267;
    end
 end
 assign n_1268 = cadence_register_n_1268;
reg cadence_register_n_1269;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1269 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1269 <= T_12_0_;
    end
 end
 assign n_1269 = cadence_register_n_1269;
reg cadence_register_n_1270;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1270 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1270 <= n_1269;
    end
 end
 assign n_1270 = cadence_register_n_1270;
reg cadence_register_n_1271;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1271 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1271 <= n_1270;
    end
 end
 assign n_1271 = cadence_register_n_1271;
reg cadence_register_n_1272;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1272 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1272 <= in1[31];
    end
 end
 assign n_1272 = cadence_register_n_1272;
reg cadence_register_n_1273;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1273 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1273 <= n_1272;
    end
 end
 assign n_1273 = cadence_register_n_1273;
reg cadence_register_n_1274;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1274 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1274 <= n_1273;
    end
 end
 assign n_1274 = cadence_register_n_1274;
reg cadence_register_n_1275;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1275 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1275 <= n_1274;
    end
 end
 assign n_1275 = cadence_register_n_1275;
reg cadence_register_n_1276;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1276 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1276 <= n_1275;
    end
 end
 assign n_1276 = cadence_register_n_1276;
reg cadence_register_n_1277;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1277 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1277 <= sub_1160_30_n_56;
    end
 end
 assign n_1277 = cadence_register_n_1277;
reg cadence_register_n_1278;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1278 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1278 <= n_1277;
    end
 end
 assign n_1278 = cadence_register_n_1278;
reg cadence_register_n_1279;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1279 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1279 <= n_1278;
    end
 end
 assign n_1279 = cadence_register_n_1279;
reg cadence_register_n_1280;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1280 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1280 <= n_1279;
    end
 end
 assign n_1280 = cadence_register_n_1280;
reg cadence_register_n_1281;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1281 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1281 <= n_1280;
    end
 end
 assign n_1281 = cadence_register_n_1281;
reg cadence_register_n_1282;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1282 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1282 <= T_4_0_;
    end
 end
 assign n_1282 = cadence_register_n_1282;
reg cadence_register_n_1283;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1283 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1283 <= n_1282;
    end
 end
 assign n_1283 = cadence_register_n_1283;
reg cadence_register_n_1284;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1284 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1284 <= n_1283;
    end
 end
 assign n_1284 = cadence_register_n_1284;
reg cadence_register_n_1285;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1285 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1285 <= n_1284;
    end
 end
 assign n_1285 = cadence_register_n_1285;
reg cadence_register_n_1286;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1286 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1286 <= n_1285;
    end
 end
 assign n_1286 = cadence_register_n_1286;
reg cadence_register_n_1287;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1287 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1287 <= T_10_0_;
    end
 end
 assign n_1287 = cadence_register_n_1287;
reg cadence_register_n_1288;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1288 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1288 <= n_1287;
    end
 end
 assign n_1288 = cadence_register_n_1288;
reg cadence_register_n_1289;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1289 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1289 <= n_1288;
    end
 end
 assign n_1289 = cadence_register_n_1289;
reg cadence_register_n_1290;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1290 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1290 <= T_24_3_;
    end
 end
 assign n_1290 = cadence_register_n_1290;
reg cadence_register_n_1291;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1291 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1291 <= in1[23];
    end
 end
 assign n_1291 = cadence_register_n_1291;
reg cadence_register_n_1292;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1292 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1292 <= n_1291;
    end
 end
 assign n_1292 = cadence_register_n_1292;
reg cadence_register_n_1293;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1293 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1293 <= n_1292;
    end
 end
 assign n_1293 = cadence_register_n_1293;
reg cadence_register_n_1294;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1294 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1294 <= n_1293;
    end
 end
 assign n_1294 = cadence_register_n_1294;
reg cadence_register_n_1295;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1295 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1295 <= n_1294;
    end
 end
 assign n_1295 = cadence_register_n_1295;
reg cadence_register_n_1296;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1296 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1296 <= in1[28];
    end
 end
 assign n_1296 = cadence_register_n_1296;
reg cadence_register_n_1297;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1297 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1297 <= n_1296;
    end
 end
 assign n_1297 = cadence_register_n_1297;
reg cadence_register_n_1298;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1298 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1298 <= n_1297;
    end
 end
 assign n_1298 = cadence_register_n_1298;
reg cadence_register_n_1299;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1299 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1299 <= n_1298;
    end
 end
 assign n_1299 = cadence_register_n_1299;
reg cadence_register_n_1300;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1300 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1300 <= n_1299;
    end
 end
 assign n_1300 = cadence_register_n_1300;
reg cadence_register_n_1301;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1301 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1301 <= in1[19];
    end
 end
 assign n_1301 = cadence_register_n_1301;
reg cadence_register_n_1302;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1302 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1302 <= n_1301;
    end
 end
 assign n_1302 = cadence_register_n_1302;
reg cadence_register_n_1303;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1303 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1303 <= n_1302;
    end
 end
 assign n_1303 = cadence_register_n_1303;
reg cadence_register_n_1304;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1304 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1304 <= n_1303;
    end
 end
 assign n_1304 = cadence_register_n_1304;
reg cadence_register_n_1305;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1305 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1305 <= n_1304;
    end
 end
 assign n_1305 = cadence_register_n_1305;
reg cadence_register_n_1306;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1306 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1306 <= sub_1070_33_n_65;
    end
 end
 assign n_1306 = cadence_register_n_1306;
reg cadence_register_n_1307;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1307 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1307 <= n_1306;
    end
 end
 assign n_1307 = cadence_register_n_1307;
reg cadence_register_n_1308;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1308 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1308 <= n_1307;
    end
 end
 assign n_1308 = cadence_register_n_1308;
reg cadence_register_n_1309;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1309 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1309 <= n_1308;
    end
 end
 assign n_1309 = cadence_register_n_1309;
reg cadence_register_n_1310;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1310 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1310 <= n_1309;
    end
 end
 assign n_1310 = cadence_register_n_1310;
reg cadence_register_n_1311;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1311 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1311 <= sub_710_48_n_61;
    end
 end
 assign n_1311 = cadence_register_n_1311;
reg cadence_register_n_1312;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1312 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1312 <= n_1311;
    end
 end
 assign n_1312 = cadence_register_n_1312;
reg cadence_register_n_1313;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1313 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1313 <= T_1_0_;
    end
 end
 assign n_1313 = cadence_register_n_1313;
reg cadence_register_n_1314;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1314 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1314 <= n_1313;
    end
 end
 assign n_1314 = cadence_register_n_1314;
reg cadence_register_n_1315;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1315 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1315 <= n_1314;
    end
 end
 assign n_1315 = cadence_register_n_1315;
reg cadence_register_n_1316;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1316 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1316 <= n_1315;
    end
 end
 assign n_1316 = cadence_register_n_1316;
reg cadence_register_n_1317;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1317 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1317 <= n_1316;
    end
 end
 assign n_1317 = cadence_register_n_1317;
reg cadence_register_n_1318;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1318 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1318 <= sub_650_50_n_40;
    end
 end
 assign n_1318 = cadence_register_n_1318;
reg cadence_register_n_1319;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1319 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1319 <= n_1318;
    end
 end
 assign n_1319 = cadence_register_n_1319;
reg cadence_register_n_1320;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1320 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1320 <= sub_590_52_n_28;
    end
 end
 assign n_1320 = cadence_register_n_1320;
reg cadence_register_n_1321;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1321 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1321 <= sub_560_53_n_25;
    end
 end
 assign n_1321 = cadence_register_n_1321;
reg cadence_register_n_1322;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1322 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1322 <= sub_530_54_n_24;
    end
 end
 assign n_1322 = cadence_register_n_1322;
reg cadence_register_n_1323;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1323 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1323 <= sub_500_55_n_20;
    end
 end
 assign n_1323 = cadence_register_n_1323;
reg cadence_register_n_1324;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1324 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1324 <= T_3_0_;
    end
 end
 assign n_1324 = cadence_register_n_1324;
reg cadence_register_n_1325;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1325 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1325 <= n_1324;
    end
 end
 assign n_1325 = cadence_register_n_1325;
reg cadence_register_n_1326;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1326 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1326 <= n_1325;
    end
 end
 assign n_1326 = cadence_register_n_1326;
reg cadence_register_n_1327;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1327 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1327 <= n_1326;
    end
 end
 assign n_1327 = cadence_register_n_1327;
reg cadence_register_n_1328;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1328 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1328 <= n_1327;
    end
 end
 assign n_1328 = cadence_register_n_1328;
reg cadence_register_n_1329;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1329 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1329 <= n_357;
    end
 end
 assign n_1329 = cadence_register_n_1329;
reg cadence_register_n_1330;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1330 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1330 <= n_1329;
    end
 end
 assign n_1330 = cadence_register_n_1330;
reg cadence_register_n_1331;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1331 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1331 <= n_1330;
    end
 end
 assign n_1331 = cadence_register_n_1331;
reg cadence_register_n_1332;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1332 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1332 <= n_1331;
    end
 end
 assign n_1332 = cadence_register_n_1332;
reg cadence_register_n_1333;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1333 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1333 <= n_1332;
    end
 end
 assign n_1333 = cadence_register_n_1333;
reg cadence_register_n_1334;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1334 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1334 <= in2[1];
    end
 end
 assign n_1334 = cadence_register_n_1334;
reg cadence_register_n_1335;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1335 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1335 <= n_1334;
    end
 end
 assign n_1335 = cadence_register_n_1335;
reg cadence_register_n_1336;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1336 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1336 <= n_1335;
    end
 end
 assign n_1336 = cadence_register_n_1336;
reg cadence_register_n_1337;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1337 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1337 <= n_1336;
    end
 end
 assign n_1337 = cadence_register_n_1337;
reg cadence_register_n_1338;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1338 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1338 <= n_1337;
    end
 end
 assign n_1338 = cadence_register_n_1338;
reg cadence_register_n_1339;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1339 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1339 <= in1[4];
    end
 end
 assign n_1339 = cadence_register_n_1339;
reg cadence_register_n_1340;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1340 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1340 <= n_1339;
    end
 end
 assign n_1340 = cadence_register_n_1340;
reg cadence_register_n_1341;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1341 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1341 <= n_1340;
    end
 end
 assign n_1341 = cadence_register_n_1341;
reg cadence_register_n_1342;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1342 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1342 <= n_1341;
    end
 end
 assign n_1342 = cadence_register_n_1342;
reg cadence_register_n_1343;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1343 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1343 <= n_1342;
    end
 end
 assign n_1343 = cadence_register_n_1343;
reg cadence_register_n_1344;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1344 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1344 <= in1[10];
    end
 end
 assign n_1344 = cadence_register_n_1344;
reg cadence_register_n_1345;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1345 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1345 <= n_1344;
    end
 end
 assign n_1345 = cadence_register_n_1345;
reg cadence_register_n_1346;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1346 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1346 <= n_1345;
    end
 end
 assign n_1346 = cadence_register_n_1346;
reg cadence_register_n_1347;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1347 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1347 <= n_1346;
    end
 end
 assign n_1347 = cadence_register_n_1347;
reg cadence_register_n_1348;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1348 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1348 <= n_1347;
    end
 end
 assign n_1348 = cadence_register_n_1348;
reg cadence_register_n_1349;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1349 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1349 <= in1[1];
    end
 end
 assign n_1349 = cadence_register_n_1349;
reg cadence_register_n_1350;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1350 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1350 <= n_1349;
    end
 end
 assign n_1350 = cadence_register_n_1350;
reg cadence_register_n_1351;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1351 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1351 <= n_1350;
    end
 end
 assign n_1351 = cadence_register_n_1351;
reg cadence_register_n_1352;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1352 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1352 <= n_1351;
    end
 end
 assign n_1352 = cadence_register_n_1352;
reg cadence_register_n_1353;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1353 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1353 <= n_1352;
    end
 end
 assign n_1353 = cadence_register_n_1353;
reg cadence_register_n_1354;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1354 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1354 <= sub_770_46_n_42;
    end
 end
 assign n_1354 = cadence_register_n_1354;
reg cadence_register_n_1355;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1355 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1355 <= sub_1130_31_n_53;
    end
 end
 assign n_1355 = cadence_register_n_1355;
reg cadence_register_n_1356;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1356 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1356 <= n_1355;
    end
 end
 assign n_1356 = cadence_register_n_1356;
reg cadence_register_n_1357;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1357 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1357 <= n_1356;
    end
 end
 assign n_1357 = cadence_register_n_1357;
reg cadence_register_n_1358;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1358 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1358 <= n_1357;
    end
 end
 assign n_1358 = cadence_register_n_1358;
reg cadence_register_n_1359;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1359 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1359 <= n_1358;
    end
 end
 assign n_1359 = cadence_register_n_1359;
reg cadence_register_n_1360;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1360 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1360 <= in1[29];
    end
 end
 assign n_1360 = cadence_register_n_1360;
reg cadence_register_n_1361;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1361 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1361 <= n_1360;
    end
 end
 assign n_1361 = cadence_register_n_1361;
reg cadence_register_n_1362;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1362 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1362 <= n_1361;
    end
 end
 assign n_1362 = cadence_register_n_1362;
reg cadence_register_n_1363;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1363 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1363 <= n_1362;
    end
 end
 assign n_1363 = cadence_register_n_1363;
reg cadence_register_n_1364;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1364 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1364 <= n_1363;
    end
 end
 assign n_1364 = cadence_register_n_1364;
reg cadence_register_n_1365;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1365 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1365 <= in1[21];
    end
 end
 assign n_1365 = cadence_register_n_1365;
reg cadence_register_n_1366;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1366 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1366 <= n_1365;
    end
 end
 assign n_1366 = cadence_register_n_1366;
reg cadence_register_n_1367;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1367 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1367 <= n_1366;
    end
 end
 assign n_1367 = cadence_register_n_1367;
reg cadence_register_n_1368;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1368 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1368 <= n_1367;
    end
 end
 assign n_1368 = cadence_register_n_1368;
reg cadence_register_n_1369;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1369 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1369 <= n_1368;
    end
 end
 assign n_1369 = cadence_register_n_1369;
reg cadence_register_n_1370;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1370 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1370 <= in1[25];
    end
 end
 assign n_1370 = cadence_register_n_1370;
reg cadence_register_n_1371;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1371 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1371 <= n_1370;
    end
 end
 assign n_1371 = cadence_register_n_1371;
reg cadence_register_n_1372;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1372 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1372 <= n_1371;
    end
 end
 assign n_1372 = cadence_register_n_1372;
reg cadence_register_n_1373;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1373 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1373 <= n_1372;
    end
 end
 assign n_1373 = cadence_register_n_1373;
reg cadence_register_n_1374;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1374 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1374 <= n_1373;
    end
 end
 assign n_1374 = cadence_register_n_1374;
reg cadence_register_n_1375;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1375 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1375 <= T_9_0_;
    end
 end
 assign n_1375 = cadence_register_n_1375;
reg cadence_register_n_1376;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1376 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1376 <= n_1375;
    end
 end
 assign n_1376 = cadence_register_n_1376;
reg cadence_register_n_1377;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1377 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1377 <= n_1376;
    end
 end
 assign n_1377 = cadence_register_n_1377;
reg cadence_register_n_1378;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1378 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1378 <= n_1377;
    end
 end
 assign n_1378 = cadence_register_n_1378;
reg cadence_register_n_1379;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1379 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1379 <= T_2_0_;
    end
 end
 assign n_1379 = cadence_register_n_1379;
reg cadence_register_n_1380;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1380 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1380 <= n_1379;
    end
 end
 assign n_1380 = cadence_register_n_1380;
reg cadence_register_n_1381;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1381 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1381 <= n_1380;
    end
 end
 assign n_1381 = cadence_register_n_1381;
reg cadence_register_n_1382;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1382 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1382 <= n_1381;
    end
 end
 assign n_1382 = cadence_register_n_1382;
reg cadence_register_n_1383;
 always @(posedge clk or negedge clr) begin
    if (clr == 1'B0) begin
       cadence_register_n_1383 <= 1'B0;
    end
    else begin
       if (stall == 1'B0) 
          cadence_register_n_1383 <= n_1382;
    end
 end
 assign n_1383 = cadence_register_n_1383;
 assign Q_0_ = ~T_0_32_;
 assign R_7_9_ = ~(n_713 & (~T_7_9_ | n_692));
 assign R_7_21_ = ~(n_711 & ~n_716);
 assign R_7_18_ = ~(n_718 & (T_7_32_ | n_693));
 assign R_7_11_ = ~(n_717 & (~T_7_11_ | n_692));
 assign R_7_17_ = ~(n_714 & (T_7_32_ | n_694));
 assign R_7_10_ = ~(n_720 & (~T_7_10_ | n_692));
 assign R_7_16_ = ~(n_712 & (~T_7_16_ | n_692));
 assign R_7_8_ = ~(n_710 & (~T_7_8_ | n_692));
 assign R_7_7_ = ~(n_685 & ~(R_8_6_ & T_7_32_));
 assign R_7_15_ = ~(n_706 & ~n_708);
 assign R_7_23_ = ~(n_687 & ~n_686);
 assign R_7_22_ = ~(n_701 & ~n_691);
 assign R_7_19_ = ~(n_698 & ~n_690);
 assign R_7_3_ = ~(n_688 & (~T_7_3_ | T_7_32_));
 assign R_7_1_ = ~(n_699 & (~T_7_1_ | T_7_32_));
 assign R_7_12_ = ~(n_702 & (~T_7_12_ | n_692));
 assign n_720 = ~(R_8_9_ & T_7_32_);
 assign n_719 = ~(R_8_23_ & n_696);
 assign n_718 = ~(R_8_17_ & T_7_32_);
 assign n_717 = ~(R_8_10_ & T_7_32_);
 assign n_716 = ~(n_695 | ~R_8_20_);
 assign n_715 = ~(R_8_3_ & T_7_32_);
 assign n_714 = ~(R_8_16_ & T_7_32_);
 assign n_713 = ~(R_8_8_ & T_7_32_);
 assign n_712 = ~(R_8_15_ & n_692);
 assign n_711 = ~(n_697 & T_7_21_);
 assign n_710 = ~(R_8_7_ & T_7_32_);
 assign n_709 = ~(R_8_19_ & n_692);
 assign n_708 = ~(n_695 | ~R_8_14_);
 assign n_707 = ~(R_8_4_ & T_7_32_);
 assign n_706 = ~(n_697 & T_7_15_);
 assign n_705 = ~(R_8_1_ & T_7_32_);
 assign n_704 = ~(R_8_13_ & T_7_32_);
 assign n_703 = ~(R_8_5_ & T_7_32_);
 assign n_702 = ~(R_8_11_ & T_7_32_);
 assign n_701 = ~(T_7_22_ & ~T_7_32_);
 assign n_700 = ~(R_8_12_ & T_7_32_);
 assign n_699 = ~(R_8_0_ & T_7_32_);
 assign n_698 = ~(T_7_19_ & ~T_7_32_);
 assign n_696 = ~n_697;
 assign n_697 = ~T_7_32_;
 assign n_692 = ~n_695;
 assign n_695 = ~T_7_32_;
 assign n_694 = ~T_7_17_;
 assign n_693 = ~T_7_18_;
 assign n_691 = (R_8_21_ & T_7_32_);
 assign n_690 = (R_8_18_ & T_7_32_);
 assign R_7_14_ = ~(n_704 & (~T_7_14_ | T_7_32_));
 assign R_7_13_ = ~(n_700 & (~T_7_13_ | T_7_32_));
 assign R_7_6_ = ~(n_703 & (~T_7_6_ | T_7_32_));
 assign n_689 = ~(T_7_32_ & n_1143);
 assign R_7_24_ = ~(n_719 & (~T_7_24_ | n_696));
 assign R_7_20_ = ~(n_709 & (~T_7_20_ | n_696));
 assign n_688 = ~(T_7_32_ & R_8_2_);
 assign n_687 = ~(T_7_23_ & ~n_696);
 assign R_7_4_ = ~(n_715 & (~T_7_4_ | T_7_32_));
 assign R_7_0_ = ~(n_689 & (~n_1160 | T_7_32_));
 assign n_686 = ~(n_697 | ~R_8_22_);
 assign R_7_5_ = ~(n_707 & (~T_7_5_ | T_7_32_));
 assign R_7_2_ = ~(n_705 & (~T_7_2_ | T_7_32_));
 assign n_685 = ~(n_695 & T_7_7_);
 assign R_8_8_ = ~(n_656 & n_678);
 assign R_8_20_ = ~(n_677 & (n_661 | n_659));
 assign R_8_16_ = ~(n_648 & ~(R_9_15_ & T_8_32_));
 assign R_8_23_ = ~(n_684 & ~n_649);
 assign R_8_19_ = ~(n_672 & ~n_652);
 assign R_8_15_ = ~(n_674 & n_679);
 assign R_8_6_ = ~(n_654 & n_673);
 assign R_8_14_ = ~(n_671 & (T_8_32_ | n_660));
 assign R_8_13_ = ~(n_669 & (T_8_32_ | n_658));
 assign R_8_21_ = ~(n_665 & ~n_655);
 assign R_8_4_ = ~(n_651 & n_670);
 assign R_8_18_ = ~(n_664 & (T_8_32_ | n_657));
 assign R_8_12_ = ~(n_650 & n_663);
 assign R_8_0_ = ~(n_653 & (~n_1203 | T_8_32_));
 assign n_684 = ~(n_659 & T_8_23_);
 assign n_683 = ~(R_9_21_ & T_8_32_);
 assign n_682 = ~(R_9_16_ & T_8_32_);
 assign n_681 = ~(R_9_9_ & T_8_32_);
 assign n_680 = ~(R_9_8_ & T_8_32_);
 assign n_679 = ~(R_9_14_ & T_8_32_);
 assign n_678 = ~(R_9_7_ & T_8_32_);
 assign n_677 = ~(n_659 & T_8_20_);
 assign n_676 = ~(R_9_6_ & T_8_32_);
 assign n_675 = ~(R_9_0_ & T_8_32_);
 assign n_674 = ~(n_659 & T_8_15_);
 assign n_673 = ~(R_9_5_ & T_8_32_);
 assign n_672 = ~(T_8_19_ & ~T_8_32_);
 assign n_671 = ~(R_9_13_ & T_8_32_);
 assign n_670 = ~(R_9_3_ & T_8_32_);
 assign n_669 = ~(R_9_12_ & T_8_32_);
 assign n_668 = ~(R_9_10_ & T_8_32_);
 assign n_667 = ~(R_9_1_ & T_8_32_);
 assign n_666 = ~(R_9_2_ & T_8_32_);
 assign n_665 = ~(n_659 & T_8_21_);
 assign n_664 = ~(R_9_17_ & T_8_32_);
 assign n_663 = ~(R_9_11_ & T_8_32_);
 assign n_662 = ~(R_9_4_ & T_8_32_);
 assign n_661 = ~R_9_19_;
 assign n_660 = ~T_8_14_;
 assign n_659 = ~T_8_32_;
 assign n_658 = ~T_8_13_;
 assign n_657 = ~T_8_18_;
 assign R_8_10_ = ~(n_681 & (~T_8_10_ | T_8_32_));
 assign R_8_17_ = ~(n_682 & (~T_8_17_ | T_8_32_));
 assign n_656 = ~(n_659 & T_8_8_);
 assign R_8_1_ = ~(n_675 & (~T_8_1_ | T_8_32_));
 assign R_8_7_ = ~(n_676 & (~T_8_7_ | T_8_32_));
 assign n_655 = ~(n_659 | ~R_9_20_);
 assign n_654 = ~(n_659 & T_8_6_);
 assign n_653 = ~(T_8_32_ & n_1195);
 assign n_652 = ~(n_659 | ~R_9_18_);
 assign R_8_2_ = ~(n_667 & (~T_8_2_ | T_8_32_));
 assign R_8_11_ = ~(n_668 & (~T_8_11_ | T_8_32_));
 assign n_651 = ~(n_659 & T_8_4_);
 assign n_650 = ~(n_659 & T_8_12_);
 assign n_649 = ~(n_659 | ~R_9_22_);
 assign R_8_9_ = ~(n_680 & (~T_8_9_ | T_8_32_));
 assign R_8_22_ = ~(n_683 & (~T_8_22_ | T_8_32_));
 assign R_8_5_ = ~(n_662 & (~T_8_5_ | T_8_32_));
 assign n_648 = ~(n_659 & T_8_16_);
 assign R_8_3_ = ~(n_666 & (~T_8_3_ | T_8_32_));
 assign R_6_25_ = ~(n_633 & ~n_641);
 assign R_6_19_ = ~(n_643 & ~n_644);
 assign R_6_12_ = ~(n_642 & (~T_6_12_ | n_622));
 assign R_6_11_ = ~(n_640 & (~T_6_11_ | n_622));
 assign R_6_10_ = ~(n_638 & (~T_6_10_ | n_622));
 assign R_6_21_ = ~(n_630 & ~n_631);
 assign R_6_9_ = ~(n_636 & (~T_6_9_ | n_622));
 assign R_6_7_ = ~(n_632 & (~T_6_7_ | n_618));
 assign R_6_23_ = ~(n_626 & ~n_617);
 assign R_6_15_ = ~(n_627 & ~n_615);
 assign R_6_14_ = ~(n_612 & (n_618 | n_623));
 assign R_6_13_ = ~(n_637 & (~T_6_13_ | n_622));
 assign n_647 = ~(R_7_21_ & n_622);
 assign n_646 = ~(R_7_4_ & T_6_32_);
 assign n_645 = ~(R_7_23_ & n_618);
 assign n_644 = ~(n_620 | ~R_7_18_);
 assign n_643 = ~(n_619 & T_6_19_);
 assign n_642 = ~(R_7_11_ & n_618);
 assign n_641 = ~(n_620 | ~R_7_24_);
 assign n_640 = ~(R_7_10_ & n_618);
 assign n_639 = ~(R_7_17_ & n_618);
 assign n_638 = ~(R_7_9_ & n_618);
 assign n_637 = ~(R_7_12_ & n_618);
 assign n_636 = ~(R_7_8_ & T_6_32_);
 assign n_635 = ~(R_7_16_ & n_618);
 assign n_634 = ~(R_7_1_ & T_6_32_);
 assign n_633 = ~(n_619 & T_6_25_);
 assign n_632 = ~(R_7_6_ & T_6_32_);
 assign n_631 = ~(n_620 | ~R_7_20_);
 assign n_630 = ~(n_619 & T_6_21_);
 assign n_629 = ~(R_7_5_ & T_6_32_);
 assign n_628 = ~(R_7_3_ & T_6_32_);
 assign n_627 = ~(n_620 & T_6_15_);
 assign n_626 = ~(T_6_23_ & ~n_622);
 assign n_625 = ~(R_7_19_ & n_622);
 assign n_624 = ~(R_7_7_ & T_6_32_);
 assign n_623 = ~T_6_14_;
 assign n_622 = ~n_621;
 assign n_621 = ~T_6_32_;
 assign n_618 = ~n_619;
 assign n_619 = ~T_6_32_;
 assign n_620 = ~T_6_32_;
 assign R_6_1_ = ~(n_611 & (~T_6_1_ | T_6_32_));
 assign R_6_3_ = ~(n_613 & (~T_6_3_ | T_6_32_));
 assign n_617 = ~(n_620 | ~R_7_22_);
 assign R_6_18_ = ~(n_639 & (~T_6_18_ | n_622));
 assign R_6_22_ = ~(n_647 & (~T_6_22_ | n_622));
 assign R_6_8_ = ~(n_624 & (~T_6_8_ | T_6_32_));
 assign n_616 = ~(T_6_32_ & n_1224);
 assign R_6_16_ = ~(n_614 & (~T_6_16_ | T_6_32_));
 assign R_6_5_ = ~(n_646 & (~T_6_5_ | T_6_32_));
 assign R_6_2_ = ~(n_634 & (~T_6_2_ | T_6_32_));
 assign R_6_0_ = ~(n_616 & (~n_1232 | T_6_32_));
 assign n_615 = ~(n_621 | ~R_7_14_);
 assign R_6_20_ = ~(n_625 & (~T_6_20_ | n_622));
 assign R_6_17_ = ~(n_635 & (~T_6_17_ | n_622));
 assign R_6_24_ = ~(n_645 & (~T_6_24_ | n_622));
 assign n_614 = ~(T_6_32_ & R_7_15_);
 assign R_6_6_ = ~(n_629 & (~T_6_6_ | T_6_32_));
 assign n_613 = ~(T_6_32_ & R_7_2_);
 assign R_6_4_ = ~(n_628 & (~T_6_4_ | T_6_32_));
 assign n_612 = ~(T_6_32_ & R_7_13_);
 assign n_611 = ~(T_6_32_ & R_7_0_);
 assign R_9_19_ = ~(n_610 & ~n_607);
 assign R_9_15_ = ~(n_603 & ~n_576);
 assign R_9_22_ = ~(n_602 & ~n_577);
 assign R_9_18_ = ~(n_600 & (n_586 | n_582));
 assign R_9_14_ = ~(n_608 & (T_9_32_ | n_591));
 assign R_9_21_ = ~(n_594 & ~n_573);
 assign R_9_3_ = ~(n_598 & n_599);
 assign R_9_13_ = ~(n_578 & ~(n_944 & T_9_32_));
 assign R_9_12_ = ~(n_580 & ~(n_940 & T_9_32_));
 assign R_9_1_ = ~(n_604 & n_595);
 assign R_9_11_ = ~((n_942 | n_585) & (T_9_32_ | n_583));
 assign n_610 = ~(n_585 & T_9_19_);
 assign n_609 = ~(n_924 & T_9_32_);
 assign n_608 = ~(n_955 & T_9_32_);
 assign n_607 = ~(n_587 | ~n_918);
 assign n_606 = ~(n_934 & T_9_32_);
 assign n_605 = ~(n_960 & T_9_32_);
 assign n_604 = ~(n_588 & ~n_950);
 assign n_603 = ~(n_585 & T_9_15_);
 assign n_602 = ~(n_585 & T_9_22_);
 assign n_601 = ~(n_954 & T_9_32_);
 assign n_600 = ~(n_907 & n_584);
 assign n_599 = ~(n_953 & T_9_32_);
 assign n_598 = ~(n_585 & ~n_951);
 assign n_597 = ~(T_9_32_ & ~n_964);
 assign n_596 = ~(n_923 & n_586);
 assign n_595 = ~(n_948 & T_9_32_);
 assign n_594 = ~(n_585 & T_9_21_);
 assign n_593 = ~R_10_1_;
 assign n_592 = ~T_9_1_;
 assign n_591 = ~T_9_14_;
 assign n_590 = ~T_9_3_;
 assign n_589 = ~R_10_10_;
 assign n_588 = ~T_9_32_;
 assign n_586 = ~n_587;
 assign n_587 = ~T_9_32_;
 assign n_584 = ~n_585;
 assign n_585 = ~T_9_32_;
 assign n_583 = ~T_9_11_;
 assign n_582 = ~T_9_18_;
 assign R_9_17_ = ~(n_575 & (~T_9_17_ | n_584));
 assign R_9_9_ = ~(n_609 & (~n_929 | T_9_32_));
 assign R_9_16_ = ~(n_571 & (~T_9_16_ | T_9_32_));
 assign n_581 = ~(T_9_32_ & n_943);
 assign n_580 = ~(n_926 & ~T_9_32_);
 assign n_579 = ~(T_9_32_ & n_1237);
 assign R_9_5_ = ~(n_572 & (~n_935 | T_9_32_));
 assign n_578 = ~(T_9_13_ & ~T_9_32_);
 assign R_9_20_ = ~(n_596 & (~T_9_20_ | n_586));
 assign R_9_4_ = ~(n_601 & (~n_952 | T_9_32_));
 assign n_577 = ~(n_587 | ~n_917);
 assign R_9_0_ = ~(n_579 & (~n_1378 | T_9_32_));
 assign R_9_8_ = ~(n_606 & (~n_912 | T_9_32_));
 assign n_576 = ~(n_587 | ~n_921);
 assign R_9_6_ = ~(n_605 & (~n_933 | T_9_32_));
 assign n_575 = ~(n_584 & n_945);
 assign n_574 = ~(T_9_32_ & n_930);
 assign n_573 = ~(n_587 | ~n_936);
 assign n_572 = ~(T_9_32_ & n_910);
 assign R_9_10_ = ~(n_574 & (~n_931 | T_9_32_));
 assign n_571 = ~(T_9_32_ & n_938);
 assign R_9_7_ = ~(n_581 & (~n_911 | T_9_32_));
 assign R_9_2_ = ~(n_597 & (~n_949 | T_9_32_));
 assign R_5_26_ = ~(n_557 & ~n_569);
 assign R_5_23_ = ~(n_560 & ~(R_6_22_ & n_535));
 assign R_5_13_ = ~(n_566 & (~T_5_13_ | n_533));
 assign R_5_0_ = ~(n_565 & n_520);
 assign R_5_19_ = ~(n_561 & ~n_563);
 assign R_5_12_ = ~(n_518 & n_564);
 assign R_5_22_ = ~(n_517 & (n_532 | n_528));
 assign R_5_10_ = ~(n_523 & (~T_5_10_ | n_533));
 assign R_5_9_ = ~(n_522 & n_542);
 assign R_5_25_ = ~(n_559 & ~n_516);
 assign R_5_24_ = ~(n_550 & (n_535 | n_541));
 assign R_5_7_ = ~(n_553 & (~T_5_7_ | n_535));
 assign R_5_6_ = ~(n_552 & n_567);
 assign R_5_21_ = ~(n_545 & ~n_548);
 assign R_5_16_ = ~(n_525 & n_551);
 assign R_5_5_ = ~(n_519 & n_549);
 assign R_5_15_ = ~(n_543 & ~n_544);
 assign R_5_4_ = ~(n_546 & n_547);
 assign R_5_3_ = ~(n_526 & ~(R_6_2_ & T_5_32_));
 assign R_5_2_ = ~(n_524 & n_555);
 assign R_5_8_ = ~(n_515 & n_556);
 assign n_570 = ~(R_6_0_ & T_5_32_);
 assign n_569 = ~(n_530 | ~R_6_25_);
 assign n_568 = ~(R_6_19_ & n_539);
 assign n_567 = ~(R_6_5_ & T_5_32_);
 assign n_566 = ~(R_6_12_ & n_539);
 assign n_565 = ~(n_538 & ~n_1047);
 assign n_564 = ~(R_6_11_ & n_532);
 assign n_563 = ~(n_537 | ~R_6_18_);
 assign n_562 = ~(R_6_10_ & T_5_32_);
 assign n_561 = ~(n_537 & T_5_19_);
 assign n_560 = ~(n_530 & T_5_23_);
 assign n_559 = ~(T_5_25_ & ~n_535);
 assign n_558 = ~(n_534 & T_5_18_);
 assign n_557 = ~(n_530 & T_5_26_);
 assign n_556 = ~(R_6_7_ & n_532);
 assign n_555 = ~(R_6_1_ & T_5_32_);
 assign n_554 = ~(R_6_16_ & n_539);
 assign n_553 = ~(R_6_6_ & n_532);
 assign n_552 = ~(n_534 & ~n_540);
 assign n_551 = ~(R_6_15_ & n_532);
 assign n_550 = ~(R_6_23_ & n_533);
 assign n_549 = ~(R_6_4_ & T_5_32_);
 assign n_548 = ~(n_537 | ~R_6_20_);
 assign n_547 = ~(R_6_3_ & n_539);
 assign n_546 = ~(n_534 & ~n_527);
 assign n_545 = ~(n_530 & T_5_21_);
 assign n_544 = ~(n_536 | ~R_6_14_);
 assign n_543 = ~(n_537 & T_5_15_);
 assign n_542 = ~(R_6_8_ & n_532);
 assign n_541 = ~T_5_24_;
 assign n_540 = ~T_5_6_;
 assign n_539 = ~n_538;
 assign n_538 = ~T_5_32_;
 assign n_537 = ~T_5_32_;
 assign n_535 = ~n_536;
 assign n_536 = ~T_5_32_;
 assign n_533 = ~n_534;
 assign n_534 = ~T_5_32_;
 assign n_532 = ~n_531;
 assign n_530 = ~n_532;
 assign n_531 = ~T_5_32_;
 assign n_529 = ~T_5_0_;
 assign n_528 = ~T_5_22_;
 assign n_527 = ~T_5_4_;
 assign R_5_20_ = ~(n_568 & (~T_5_20_ | n_532));
 assign R_5_17_ = ~(n_554 & (~T_5_17_ | n_533));
 assign n_526 = ~(n_538 & T_5_3_);
 assign n_525 = ~(n_534 & T_5_16_);
 assign n_524 = ~(n_531 & T_5_2_);
 assign n_523 = ~(n_532 & R_6_9_);
 assign n_522 = ~(n_536 & T_5_9_);
 assign n_521 = ~(T_5_32_ & R_6_13_);
 assign n_520 = ~(T_5_32_ & n_1038);
 assign R_5_14_ = ~(n_521 & (~T_5_14_ | n_539));
 assign n_519 = ~(n_536 & T_5_5_);
 assign n_518 = ~(n_536 & T_5_12_);
 assign n_517 = ~(n_539 & R_6_21_);
 assign n_516 = ~(n_530 | ~R_6_24_);
 assign R_5_11_ = ~(n_562 & (~T_5_11_ | n_532));
 assign R_5_18_ = ~(n_558 & (~R_6_17_ | n_537));
 assign n_515 = ~(n_537 & T_5_8_);
 assign R_5_1_ = ~(n_570 & (~T_5_1_ | T_5_32_));
 assign R_10_7_ = ~(n_510 & (~T_10_7_ | n_490));
 assign R_10_15_ = ~(n_512 & ~n_514);
 assign R_10_8_ = ~(n_482 & ~(R_11_7_ & n_492));
 assign R_10_14_ = ~((n_485 | n_489) & (n_493 | n_498));
 assign R_10_21_ = ~(n_502 & ~n_481);
 assign R_10_13_ = ~(n_513 & (n_493 | n_486));
 assign R_10_4_ = ~((n_496 | n_489) & (T_10_32_ | n_487));
 assign R_10_20_ = ((R_11_19_ & n_490) | ~(n_493 | n_495));
 assign R_10_19_ = ~(n_501 & ~n_479);
 assign R_10_11_ = ~((n_488 | n_489) & (n_490 | n_494));
 assign R_10_0_ = ~(n_483 & (~n_1289 | T_10_32_));
 assign R_10_9_ = ~(n_478 & n_504);
 assign n_514 = ~(n_497 | n_489);
 assign n_513 = ~(R_11_12_ & n_492);
 assign n_512 = ~(n_489 & T_10_15_);
 assign n_511 = ~(R_11_17_ & n_493);
 assign n_510 = ~(R_11_6_ & n_492);
 assign n_509 = ~(R_11_5_ & n_490);
 assign n_508 = ~(R_11_0_ & T_10_32_);
 assign n_507 = ~(R_11_1_ & T_10_32_);
 assign n_506 = ~(R_11_2_ & T_10_32_);
 assign n_505 = ~(R_11_16_ & n_490);
 assign n_504 = ~(R_11_8_ & n_492);
 assign n_503 = ~(R_11_11_ & n_492);
 assign n_502 = ~(n_484 & T_10_21_);
 assign n_501 = ~(n_484 & T_10_19_);
 assign n_500 = ~(R_11_15_ & T_10_32_);
 assign n_499 = ~(R_11_9_ & n_492);
 assign n_498 = ~T_10_14_;
 assign n_497 = ~R_11_14_;
 assign n_496 = ~R_11_3_;
 assign n_495 = ~T_10_20_;
 assign n_494 = ~T_10_11_;
 assign n_493 = ~n_484;
 assign n_484 = ~T_10_32_;
 assign n_492 = ~n_491;
 assign n_491 = ~T_10_32_;
 assign n_490 = ~n_489;
 assign n_489 = ~T_10_32_;
 assign n_488 = ~R_11_10_;
 assign n_487 = ~T_10_4_;
 assign n_486 = ~T_10_13_;
 assign n_485 = ~R_11_13_;
 assign n_483 = ~(T_10_32_ & n_1206);
 assign n_482 = ~(n_484 & T_10_8_);
 assign R_10_1_ = ~(n_508 & (~T_10_1_ | T_10_32_));
 assign R_10_12_ = ~(n_503 & (~T_10_12_ | n_490));
 assign R_10_6_ = ~(n_509 & (~T_10_6_ | n_490));
 assign R_10_18_ = ~(n_511 & (~T_10_18_ | n_493));
 assign R_10_2_ = ~(n_507 & (~T_10_2_ | T_10_32_));
 assign R_10_10_ = ~(n_499 & (~T_10_10_ | n_492));
 assign R_10_3_ = ~(n_506 & (~T_10_3_ | T_10_32_));
 assign n_481 = ~(n_489 | ~R_11_20_);
 assign R_10_17_ = ~(n_505 & (~T_10_17_ | n_493));
 assign n_480 = ~(T_10_32_ & R_11_4_);
 assign n_479 = ~(n_489 | ~R_11_18_);
 assign n_478 = ~(n_484 & T_10_9_);
 assign R_10_5_ = ~(n_480 & (~T_10_5_ | T_10_32_));
 assign R_10_16_ = ~(n_500 & (~T_10_16_ | n_490));
 assign R_4_24_ = ~((n_444 | n_438) & (n_435 | n_447));
 assign R_4_21_ = ~(n_475 & ~n_430);
 assign R_4_14_ = ~(n_474 & (n_440 | n_443));
 assign R_4_20_ = ~(n_471 & (n_435 | n_442));
 assign R_4_12_ = ~(n_469 & ~(n_889 & T_4_32_));
 assign R_4_23_ = ~(n_459 & ~n_462);
 assign R_4_19_ = ~(n_466 & ~n_426);
 assign R_4_10_ = ~(n_465 & (T_4_32_ | n_446));
 assign R_4_27_ = ~(n_464 & ~n_476);
 assign R_4_26_ = ~(n_467 & ~n_433);
 assign R_4_25_ = ~(n_456 & ~n_428);
 assign R_4_7_ = ~(n_424 & n_473);
 assign R_4_6_ = ~(n_434 & (T_4_32_ | n_448));
 assign R_4_16_ = ~(n_453 & (T_4_32_ | n_450));
 assign R_4_5_ = ~(n_432 & n_454);
 assign R_4_4_ = ~(n_429 & n_452);
 assign R_4_15_ = ~(n_472 & n_460);
 assign R_4_3_ = ~(n_451 & n_461);
 assign R_4_9_ = ~(n_431 & n_463);
 assign n_477 = ~(n_861 & T_4_32_);
 assign n_476 = ~(n_436 | ~n_870);
 assign n_475 = ~(n_436 & T_4_21_);
 assign n_474 = ~(n_862 & T_4_32_);
 assign n_473 = ~(n_880 & T_4_32_);
 assign n_472 = ~(T_4_15_ & ~n_435);
 assign n_471 = ~(n_854 & T_4_32_);
 assign n_470 = ~(n_901 & T_4_32_);
 assign n_469 = ~(n_436 & ~n_449);
 assign n_468 = ~(n_890 & T_4_32_);
 assign n_467 = ~(n_437 & T_4_26_);
 assign n_466 = ~(n_436 & T_4_19_);
 assign n_465 = ~(n_838 & T_4_32_);
 assign n_464 = ~(n_436 & T_4_27_);
 assign n_463 = ~(n_841 & T_4_32_);
 assign n_462 = ~(n_437 | ~n_867);
 assign n_461 = ~(n_894 & T_4_32_);
 assign n_460 = ~(n_842 & n_439);
 assign n_459 = ~(n_436 & T_4_23_);
 assign n_458 = ~(n_846 & n_435);
 assign n_457 = ~(n_849 & n_435);
 assign n_456 = ~(n_437 & T_4_25_);
 assign n_455 = ~(n_856 & n_435);
 assign n_454 = ~(n_883 & T_4_32_);
 assign n_453 = ~(n_853 & T_4_32_);
 assign n_452 = ~(n_898 & T_4_32_);
 assign n_451 = ~(n_441 & ~n_445);
 assign n_450 = ~T_4_16_;
 assign n_449 = ~T_4_12_;
 assign n_448 = ~T_4_6_;
 assign n_447 = ~T_4_24_;
 assign n_446 = ~T_4_10_;
 assign n_445 = ~n_895;
 assign n_444 = ~n_871;
 assign n_443 = ~T_4_14_;
 assign n_442 = ~T_4_20_;
 assign n_441 = ~T_4_32_;
 assign n_440 = ~n_437;
 assign n_437 = ~T_4_32_;
 assign n_439 = ~n_438;
 assign n_438 = ~T_4_32_;
 assign n_435 = ~n_436;
 assign n_436 = ~T_4_32_;
 assign R_4_1_ = ~(n_470 & (~n_902 | T_4_32_));
 assign n_434 = ~(T_4_32_ & n_879);
 assign n_433 = ~(n_438 | ~n_875);
 assign R_4_22_ = ~(n_455 & (~T_4_22_ | n_439));
 assign n_432 = ~(n_441 & T_4_5_);
 assign R_4_11_ = ~(n_468 & ~(n_437 & T_4_11_));
 assign R_4_2_ = ~(n_425 & (~n_903 | T_4_32_));
 assign n_431 = ~(n_436 & T_4_9_);
 assign R_4_18_ = ~(n_458 & (~T_4_18_ | n_439));
 assign n_430 = ~(n_438 | ~n_873);
 assign R_4_0_ = ~(n_427 & (~n_1286 | T_4_32_));
 assign n_429 = ~(n_441 & T_4_4_);
 assign n_428 = ~(n_438 | ~n_855);
 assign R_4_17_ = ~(n_457 & (~T_4_17_ | n_439));
 assign n_427 = ~(T_4_32_ & n_1126);
 assign R_4_13_ = ~(n_477 & (~T_4_13_ | n_440));
 assign n_426 = ~(n_437 | ~n_843);
 assign R_4_8_ = ~(n_423 & (~T_4_8_ | T_4_32_));
 assign n_425 = ~(T_4_32_ & n_836);
 assign n_424 = ~(n_436 & T_4_7_);
 assign n_423 = ~(T_4_32_ & n_872);
 assign R_11_14_ = ~(n_420 & (T_11_32_ | n_404));
 assign R_11_7_ = ~(n_419 & (~T_11_7_ | T_11_32_));
 assign R_11_6_ = ~(n_417 & (~T_11_6_ | T_11_32_));
 assign R_11_16_ = ~(n_400 & n_409);
 assign R_11_12_ = ~(n_396 & n_418);
 assign R_11_4_ = ~(n_414 & (~T_11_4_ | T_11_32_));
 assign R_11_11_ = ~(n_408 & (T_11_32_ | n_403));
 assign R_11_19_ = ~(n_413 & ~n_395);
 assign R_11_15_ = ~(n_405 & ~n_401);
 assign R_11_9_ = ~(n_398 & (~T_11_9_ | T_11_32_));
 assign n_422 = ~(R_12_16_ & T_11_32_);
 assign n_421 = ~(R_12_19_ & T_11_32_);
 assign n_420 = ~(R_12_13_ & T_11_32_);
 assign n_419 = ~(R_12_6_ & T_11_32_);
 assign n_418 = ~(R_12_11_ & T_11_32_);
 assign n_417 = ~(R_12_5_ & T_11_32_);
 assign n_416 = ~(R_12_12_ & T_11_32_);
 assign n_415 = ~(R_12_4_ & T_11_32_);
 assign n_414 = ~(R_12_3_ & T_11_32_);
 assign n_413 = ~(n_402 & T_11_19_);
 assign n_412 = ~(R_12_2_ & T_11_32_);
 assign n_411 = ~(R_12_7_ & T_11_32_);
 assign n_410 = ~(R_12_1_ & T_11_32_);
 assign n_409 = ~(R_12_15_ & T_11_32_);
 assign n_408 = ~(R_12_10_ & T_11_32_);
 assign n_407 = ~(R_12_0_ & T_11_32_);
 assign n_406 = ~(R_12_9_ & T_11_32_);
 assign n_405 = ~(T_11_15_ & ~T_11_32_);
 assign n_404 = ~T_11_14_;
 assign n_403 = ~T_11_11_;
 assign n_402 = ~T_11_32_;
 assign n_401 = (R_12_14_ & T_11_32_);
 assign R_11_1_ = ~(n_407 & (~T_11_1_ | T_11_32_));
 assign R_11_20_ = ~(n_421 & (~T_11_20_ | T_11_32_));
 assign n_400 = ~(n_402 & T_11_16_);
 assign n_399 = ~(T_11_32_ & n_1071);
 assign R_11_3_ = ~(n_412 & (~T_11_3_ | T_11_32_));
 assign n_398 = ~(T_11_32_ & R_12_8_);
 assign R_11_10_ = ~(n_406 & (~T_11_10_ | T_11_32_));
 assign n_397 = ~(T_11_32_ & R_12_17_);
 assign R_11_0_ = ~(n_399 & (~n_1077 | T_11_32_));
 assign R_11_13_ = ~(n_416 & (~T_11_13_ | T_11_32_));
 assign R_11_17_ = ~(n_422 & (~T_11_17_ | T_11_32_));
 assign n_396 = ~(n_402 & T_11_12_);
 assign R_11_18_ = ~(n_397 & (~T_11_18_ | T_11_32_));
 assign R_11_5_ = ~(n_415 & (~T_11_5_ | T_11_32_));
 assign R_11_8_ = ~(n_411 & (~T_11_8_ | T_11_32_));
 assign n_395 = ~(n_402 | ~R_12_18_);
 assign R_11_2_ = ~(n_410 & (~T_11_2_ | T_11_32_));
 assign R_3_25_ = ~(n_383 & ~n_355);
 assign R_3_15_ = ~(n_389 & n_391);
 assign R_3_0_ = ~(n_394 & (~n_1328 | T_3_32_));
 assign R_3_21_ = ~(n_384 & ~n_354);
 assign R_3_13_ = ~(n_385 & (T_3_32_ | n_356));
 assign R_3_12_ = ~(n_349 & n_382);
 assign R_3_28_ = ~(n_378 & ~n_348);
 assign R_3_27_ = ~(n_381 & ~n_350);
 assign R_3_8_ = ~(n_352 & n_387);
 assign R_3_23_ = ~(n_364 & ~n_353);
 assign R_3_19_ = ~(n_372 & ~n_374);
 assign R_3_7_ = ~(n_351 & n_369);
 assign R_3_17_ = ~(n_367 & (T_3_32_ | n_363));
 assign n_394 = ~(T_3_32_ & ~n_1333);
 assign n_393 = ~(R_4_2_ & T_3_32_);
 assign n_392 = ~(R_4_21_ & n_359);
 assign n_391 = ~(R_4_14_ & n_359);
 assign n_390 = ~(R_4_0_ & T_3_32_);
 assign n_389 = ~(n_362 & T_3_15_);
 assign n_388 = ~(R_4_1_ & T_3_32_);
 assign n_387 = ~(R_4_7_ & T_3_32_);
 assign n_386 = ~(R_4_13_ & T_3_32_);
 assign n_385 = ~(R_4_12_ & T_3_32_);
 assign n_384 = ~(n_362 & T_3_21_);
 assign n_383 = ~(n_362 & T_3_25_);
 assign n_382 = ~(R_4_11_ & T_3_32_);
 assign n_381 = ~(n_362 & T_3_27_);
 assign n_380 = ~(R_4_19_ & T_3_32_);
 assign n_379 = ~(R_4_10_ & T_3_32_);
 assign n_378 = ~(T_3_28_ & ~n_361);
 assign n_377 = ~(R_4_9_ & T_3_32_);
 assign n_376 = ~(R_4_15_ & T_3_32_);
 assign n_375 = ~(n_362 & T_3_24_);
 assign n_374 = ~(n_360 | ~R_4_18_);
 assign n_373 = ~(R_4_8_ & T_3_32_);
 assign n_372 = ~(T_3_19_ & ~n_361);
 assign n_371 = ~(R_4_17_ & T_3_32_);
 assign n_370 = ~(R_4_25_ & n_359);
 assign n_369 = ~(R_4_6_ & T_3_32_);
 assign n_368 = ~(R_4_5_ & T_3_32_);
 assign n_367 = ~(R_4_16_ & T_3_32_);
 assign n_366 = ~(R_4_4_ & T_3_32_);
 assign n_365 = ~(R_4_3_ & T_3_32_);
 assign n_364 = ~(T_3_23_ & ~n_361);
 assign n_363 = ~T_3_17_;
 assign n_361 = ~n_362;
 assign n_362 = ~T_3_32_;
 assign n_360 = ~T_3_32_;
 assign n_359 = ~n_358;
 assign n_358 = ~T_3_32_;
 assign n_357 = ~{in2[3]};
 assign n_356 = ~T_3_13_;
 assign R_3_4_ = ~(n_365 & (~T_3_4_ | T_3_32_));
 assign R_3_5_ = ~(n_366 & (~T_3_5_ | T_3_32_));
 assign n_355 = ~(n_360 | ~R_4_24_);
 assign n_354 = ~(n_360 | ~R_4_20_);
 assign R_3_16_ = ~(n_376 & (~T_3_16_ | n_361));
 assign n_353 = ~(n_360 | ~R_4_22_);
 assign R_3_3_ = ~(n_393 & (~T_3_3_ | T_3_32_));
 assign R_3_11_ = ~(n_379 & (~T_3_11_ | T_3_32_));
 assign R_3_20_ = ~(n_380 & (~T_3_20_ | T_3_32_));
 assign R_3_10_ = ~(n_377 & (~T_3_10_ | T_3_32_));
 assign n_352 = ~(n_362 & T_3_8_);
 assign R_3_26_ = ~(n_370 & (~T_3_26_ | n_359));
 assign R_3_18_ = ~(n_371 & (~T_3_18_ | n_361));
 assign R_3_22_ = ~(n_392 & (~T_3_22_ | n_359));
 assign R_3_1_ = ~(n_390 & (~T_3_1_ | T_3_32_));
 assign R_3_14_ = ~(n_386 & (~T_3_14_ | T_3_32_));
 assign R_3_24_ = ~(n_375 & (~R_4_23_ | n_362));
 assign n_351 = ~(n_362 & T_3_7_);
 assign R_3_6_ = ~(n_368 & (~T_3_6_ | T_3_32_));
 assign n_350 = ~(n_360 | ~R_4_26_);
 assign n_349 = ~(n_362 & T_3_12_);
 assign R_3_2_ = ~(n_388 & (~T_3_2_ | T_3_32_));
 assign R_3_9_ = ~(n_373 & (~T_3_9_ | T_3_32_));
 assign n_348 = ~(n_360 | ~R_4_27_);
 assign R_12_19_ = ~(n_336 & ~n_347);
 assign R_12_16_ = ~(n_344 & (T_12_32_ | n_318));
 assign R_12_5_ = ~(n_316 & ~(R_13_4_ & T_12_32_));
 assign R_12_15_ = ~(n_333 & ~n_334);
 assign R_12_11_ = ~(n_338 & ~(R_13_10_ & T_12_32_));
 assign R_12_3_ = ~(n_340 & n_343);
 assign R_12_18_ = ~(n_339 & ~(R_13_17_ & n_320));
 assign R_12_17_ = ~(n_330 & ~(R_13_16_ & n_320));
 assign R_12_14_ = ~(n_329 & (n_322 | n_326));
 assign R_12_8_ = ~(n_328 & (~T_12_8_ | T_12_32_));
 assign n_347 = ~(n_324 | ~R_13_18_);
 assign n_346 = ~(R_13_12_ & n_320);
 assign n_345 = ~(R_13_5_ & T_12_32_);
 assign n_344 = ~(T_12_32_ & ~n_327);
 assign n_343 = ~(R_13_2_ & T_12_32_);
 assign n_342 = ~(R_13_11_ & T_12_32_);
 assign n_341 = ~(R_13_3_ & T_12_32_);
 assign n_340 = ~(n_323 & ~n_325);
 assign n_339 = ~(n_324 & T_12_18_);
 assign n_338 = ~(n_321 & T_12_11_);
 assign n_337 = ~(R_13_9_ & T_12_32_);
 assign n_336 = ~(n_324 & T_12_19_);
 assign n_335 = ~(R_13_0_ & T_12_32_);
 assign n_334 = ~(n_324 | ~R_13_14_);
 assign n_333 = ~(T_12_15_ & ~n_322);
 assign n_332 = ~(R_13_6_ & T_12_32_);
 assign n_331 = ~(R_13_8_ & T_12_32_);
 assign n_330 = ~(n_324 & T_12_17_);
 assign n_329 = ~(R_13_13_ & n_320);
 assign n_328 = ~(R_13_7_ & T_12_32_);
 assign n_327 = ~R_13_15_;
 assign n_326 = ~T_12_14_;
 assign n_325 = ~T_12_3_;
 assign n_324 = ~T_12_32_;
 assign n_323 = ~T_12_32_;
 assign n_322 = ~n_321;
 assign n_321 = ~T_12_32_;
 assign n_320 = ~n_319;
 assign n_319 = ~T_12_32_;
 assign n_318 = ~T_12_16_;
 assign R_12_1_ = ~(n_335 & (~T_12_1_ | T_12_32_));
 assign R_12_6_ = ~(n_345 & (~T_12_6_ | n_320));
 assign n_317 = ~(T_12_32_ & n_1265);
 assign R_12_4_ = ~(n_341 & (~T_12_4_ | T_12_32_));
 assign R_12_2_ = ~(n_315 & (~T_12_2_ | T_12_32_));
 assign n_316 = ~(n_321 & T_12_5_);
 assign R_12_12_ = ~(n_342 & (~T_12_12_ | T_12_32_));
 assign R_12_10_ = ~(n_337 & (~T_12_10_ | T_12_32_));
 assign n_315 = ~(T_12_32_ & R_13_1_);
 assign R_12_0_ = ~(n_317 & (~n_1271 | T_12_32_));
 assign R_12_7_ = ~(n_332 & (~T_12_7_ | T_12_32_));
 assign R_12_9_ = ~(n_331 & (~T_12_9_ | T_12_32_));
 assign R_12_13_ = ~(n_346 & (~T_12_13_ | n_322));
 assign R_2_22_ = ~(n_301 & ~(R_3_21_ & n_276));
 assign R_2_26_ = ~(n_300 & ~n_305);
 assign R_2_23_ = ~(n_310 & ~n_311);
 assign R_2_3_ = ~(n_312 & (~T_2_3_ | T_2_32_));
 assign R_2_1_ = ~(n_272 & ~(R_3_0_ & T_2_32_));
 assign R_2_29_ = ~(n_295 & ~n_314);
 assign R_2_15_ = ~(n_304 & ~n_307);
 assign R_2_0_ = ~(n_269 & (~n_1383 | T_2_32_));
 assign R_2_25_ = ~(n_293 & ~n_271);
 assign R_2_21_ = ~(n_297 & ~(R_3_20_ & n_276));
 assign R_2_19_ = ~(n_288 & ~(R_3_18_ & n_276));
 assign R_2_28_ = ~(n_298 & ~n_313);
 assign R_2_27_ = ~(n_287 & ~n_290);
 assign R_2_10_ = ~(n_291 & (~T_2_10_ | T_2_32_));
 assign R_2_9_ = ~(n_270 & n_303);
 assign R_2_8_ = ~(n_289 & (~T_2_8_ | T_2_32_));
 assign R_2_7_ = ~(n_284 & n_285);
 assign R_2_6_ = ~(n_282 & (~T_2_6_ | T_2_32_));
 assign R_2_17_ = ~(n_280 & (n_274 | n_279));
 assign R_2_4_ = ~(n_306 & (~T_2_4_ | T_2_32_));
 assign n_314 = ~(n_273 | ~R_3_28_);
 assign n_313 = ~(n_277 | ~R_3_27_);
 assign n_312 = ~(R_3_2_ & T_2_32_);
 assign n_311 = ~(n_273 | ~R_3_22_);
 assign n_310 = ~(n_268 & T_2_23_);
 assign n_309 = ~(R_3_15_ & n_274);
 assign n_308 = ~(R_3_1_ & T_2_32_);
 assign n_307 = ~(n_277 | ~R_3_14_);
 assign n_306 = ~(R_3_3_ & T_2_32_);
 assign n_305 = ~(n_277 | ~R_3_25_);
 assign n_304 = ~(n_273 & T_2_15_);
 assign n_303 = ~(R_3_8_ & T_2_32_);
 assign n_302 = ~(R_3_13_ & T_2_32_);
 assign n_301 = ~(n_268 & T_2_22_);
 assign n_300 = ~(T_2_26_ & ~n_274);
 assign n_299 = ~(R_3_12_ & T_2_32_);
 assign n_298 = ~(T_2_28_ & ~T_2_32_);
 assign n_297 = ~(n_273 & T_2_21_);
 assign n_296 = ~(R_3_11_ & T_2_32_);
 assign n_295 = ~(n_275 & T_2_29_);
 assign n_294 = ~(R_3_10_ & T_2_32_);
 assign n_293 = ~(n_273 & T_2_25_);
 assign n_292 = ~(R_3_19_ & n_274);
 assign n_291 = ~(R_3_9_ & T_2_32_);
 assign n_290 = ~(n_273 | ~R_3_26_);
 assign n_289 = ~(R_3_7_ & T_2_32_);
 assign n_288 = ~(n_273 & T_2_19_);
 assign n_287 = ~(n_275 & T_2_27_);
 assign n_286 = ~(R_3_23_ & T_2_32_);
 assign n_285 = ~(R_3_6_ & T_2_32_);
 assign n_284 = ~(n_273 & ~n_278);
 assign n_283 = ~(R_3_17_ & n_274);
 assign n_282 = ~(R_3_5_ & T_2_32_);
 assign n_281 = ~(R_3_4_ & T_2_32_);
 assign n_280 = ~(R_3_16_ & n_274);
 assign n_279 = ~T_2_17_;
 assign n_278 = ~T_2_7_;
 assign n_277 = ~T_2_32_;
 assign n_276 = ~n_268;
 assign n_275 = ~n_276;
 assign n_268 = ~T_2_32_;
 assign n_274 = ~n_273;
 assign n_273 = ~T_2_32_;
 assign R_2_24_ = ~(n_286 & (~T_2_24_ | n_274));
 assign R_2_2_ = ~(n_308 & (~T_2_2_ | T_2_32_));
 assign R_2_14_ = ~(n_302 & (~T_2_14_ | T_2_32_));
 assign R_2_12_ = ~(n_296 & (~T_2_12_ | T_2_32_));
 assign R_2_16_ = ~(n_309 & (~T_2_16_ | n_274));
 assign n_272 = ~(T_2_1_ & ~T_2_32_);
 assign R_2_18_ = ~(n_283 & (~T_2_18_ | n_274));
 assign R_2_13_ = ~(n_299 & (~T_2_13_ | T_2_32_));
 assign n_271 = ~(n_277 | ~R_3_24_);
 assign n_270 = ~(n_273 & T_2_9_);
 assign R_2_20_ = ~(n_292 & (~T_2_20_ | n_276));
 assign R_2_11_ = ~(n_294 & (~T_2_11_ | T_2_32_));
 assign n_269 = ~(T_2_32_ & n_1250);
 assign R_2_5_ = ~(n_281 & ~(T_2_5_ & n_273));
 assign R_13_15_ = ~(n_259 & ~n_248);
 assign R_13_12_ = ~(n_265 & (~T_13_12_ | n_251));
 assign R_13_11_ = ~(n_263 & (n_251 | n_253));
 assign R_13_16_ = ~(n_255 & (~T_13_16_ | n_251));
 assign R_13_13_ = ~(n_254 & (n_251 | n_252));
 assign n_267 = ~(R_14_17_ & n_251);
 assign n_266 = ~(n_980 & n_251);
 assign n_265 = ~(R_14_11_ & T_13_32_);
 assign n_264 = ~(n_985 & T_13_32_);
 assign n_263 = ~(n_984 & T_13_32_);
 assign n_262 = ~(n_969 & T_13_32_);
 assign n_261 = ~(n_970 & T_13_32_);
 assign n_260 = ~(n_971 & T_13_32_);
 assign n_259 = ~(T_13_15_ & ~n_251);
 assign n_258 = ~(n_979 & T_13_32_);
 assign n_257 = ~(n_972 & T_13_32_);
 assign n_256 = ~(n_968 & T_13_32_);
 assign n_255 = ~(R_14_15_ & n_251);
 assign n_254 = ~(n_973 & T_13_32_);
 assign n_253 = ~T_13_11_;
 assign n_251 = ~n_250;
 assign n_250 = ~T_13_32_;
 assign n_252 = ~T_13_13_;
 assign R_13_5_ = ~(n_264 & (~T_13_5_ | T_13_32_));
 assign R_13_0_ = ~(n_249 & (~n_1156 | T_13_32_));
 assign n_249 = ~(T_13_32_ & n_1146);
 assign R_13_4_ = ~(n_245 & (~T_13_4_ | T_13_32_));
 assign n_248 = ~(n_250 | ~n_986);
 assign R_13_6_ = ~(n_260 & (~T_13_6_ | T_13_32_));
 assign R_13_17_ = ~(n_266 & (~T_13_17_ | n_251));
 assign R_13_3_ = ~(n_262 & (~T_13_3_ | T_13_32_));
 assign R_13_18_ = ~(n_267 & (~T_13_18_ | n_251));
 assign n_247 = ~(T_13_32_ & n_966);
 assign R_13_14_ = ~(n_257 & (~T_13_14_ | n_251));
 assign R_13_10_ = ~(n_261 & (~T_13_10_ | n_251));
 assign n_246 = ~(T_13_32_ & n_977);
 assign R_13_9_ = ~(n_256 & (~T_13_9_ | T_13_32_));
 assign R_13_8_ = ~(n_244 & (~T_13_8_ | T_13_32_));
 assign R_13_7_ = ~(n_246 & (~T_13_7_ | n_251));
 assign n_245 = ~(T_13_32_ & n_967);
 assign n_244 = ~(T_13_32_ & n_978);
 assign R_13_2_ = ~(n_247 & (~T_13_2_ | T_13_32_));
 assign R_13_1_ = ~(n_258 & (~T_13_1_ | T_13_32_));
 assign R_1_23_ = ~(n_232 & ~(R_2_22_ & T_1_32_));
 assign R_1_27_ = (n_243 | (n_211 & T_1_27_));
 assign R_1_30_ = ~(n_225 & ~(R_2_29_ & T_1_32_));
 assign R_1_15_ = ~(n_231 & ~(R_2_14_ & T_1_32_));
 assign R_1_26_ = ~(n_223 & ~(R_2_25_ & T_1_32_));
 assign R_1_22_ = ~(n_227 & ~(R_2_21_ & T_1_32_));
 assign R_1_14_ = ~(n_230 & (T_1_32_ | n_212));
 assign R_1_21_ = ~(n_221 & ~(R_2_20_ & T_1_32_));
 assign R_1_29_ = ~(n_229 & ~(R_2_28_ & T_1_32_));
 assign R_1_28_ = ~(n_218 & ~(R_2_27_ & T_1_32_));
 assign R_1_25_ = ~(n_228 & ~(R_2_24_ & T_1_32_));
 assign R_1_19_ = ~(n_215 & ~(R_2_18_ & T_1_32_));
 assign n_243 = ~(n_211 | ~R_2_26_);
 assign n_242 = ~(R_2_4_ & T_1_32_);
 assign n_241 = ~(R_2_3_ & T_1_32_);
 assign n_240 = ~(R_2_23_ & T_1_32_);
 assign n_239 = ~(R_2_16_ & T_1_32_);
 assign n_238 = ~(R_2_2_ & T_1_32_);
 assign n_237 = ~(T_1_32_ & n_1338);
 assign n_236 = ~(R_2_17_ & T_1_32_);
 assign n_235 = ~(R_2_15_ & T_1_32_);
 assign n_234 = ~(R_2_0_ & T_1_32_);
 assign n_233 = ~(R_2_9_ & T_1_32_);
 assign n_232 = ~(n_211 & T_1_23_);
 assign n_231 = ~(n_211 & T_1_15_);
 assign n_230 = ~(R_2_13_ & T_1_32_);
 assign n_229 = ~(n_211 & T_1_29_);
 assign n_228 = ~(n_211 & T_1_25_);
 assign n_227 = ~(n_211 & T_1_22_);
 assign n_226 = ~(R_2_12_ & T_1_32_);
 assign n_225 = ~(n_211 & T_1_30_);
 assign n_224 = ~(R_2_11_ & T_1_32_);
 assign n_223 = ~(n_211 & T_1_26_);
 assign n_222 = ~(R_2_10_ & T_1_32_);
 assign n_221 = ~(n_211 & T_1_21_);
 assign n_220 = ~(R_2_19_ & T_1_32_);
 assign n_219 = ~(R_2_8_ & T_1_32_);
 assign n_218 = ~(n_211 & T_1_28_);
 assign n_217 = ~(R_2_7_ & T_1_32_);
 assign n_216 = ~(R_2_6_ & T_1_32_);
 assign n_215 = ~(n_211 & T_1_19_);
 assign n_214 = ~(R_2_5_ & T_1_32_);
 assign n_213 = ~(R_2_1_ & T_1_32_);
 assign n_212 = ~T_1_14_;
 assign n_211 = ~T_1_32_;
 assign R_1_0_ = ~(n_237 & (~n_1317 | T_1_32_));
 assign R_1_5_ = ~(n_242 & (~T_1_5_ | T_1_32_));
 assign R_1_16_ = ~(n_235 & (~T_1_16_ | T_1_32_));
 assign R_1_18_ = ~(n_236 & (~T_1_18_ | T_1_32_));
 assign R_1_3_ = ~(n_238 & (~T_1_3_ | T_1_32_));
 assign R_1_4_ = ~(n_241 & (~T_1_4_ | T_1_32_));
 assign R_1_12_ = ~(n_224 & (~T_1_12_ | T_1_32_));
 assign R_1_2_ = ~(n_213 & (~T_1_2_ | T_1_32_));
 assign R_1_24_ = ~(n_240 & (~T_1_24_ | T_1_32_));
 assign R_1_20_ = ~(n_220 & (~T_1_20_ | T_1_32_));
 assign R_1_7_ = ~(n_216 & (~T_1_7_ | T_1_32_));
 assign R_1_1_ = ~(n_234 & (~T_1_1_ | T_1_32_));
 assign R_1_17_ = ~(n_239 & (~T_1_17_ | T_1_32_));
 assign R_1_11_ = ~(n_222 & (~T_1_11_ | T_1_32_));
 assign R_1_13_ = ~(n_226 & (~T_1_13_ | T_1_32_));
 assign R_1_9_ = ~(n_219 & (~T_1_9_ | T_1_32_));
 assign R_1_8_ = ~(n_217 & (~T_1_8_ | T_1_32_));
 assign R_1_10_ = ~(n_233 & (~T_1_10_ | T_1_32_));
 assign R_1_6_ = ~(n_214 & (~T_1_6_ | T_1_32_));
 assign Q_1_ = ~T_1_32_;
 assign Q_7_ = ~T_7_32_;
 assign Q_2_ = ~T_2_32_;
 assign Q_5_ = ~n_835;
 assign Q_4_ = ~T_4_32_;
 assign Q_3_ = ~T_3_32_;
 assign Q_6_ = ~T_6_32_;
 assign R_14_15_ = ~(n_194 & ~n_965);
 assign n_210 = ~(R_15_4_ & T_14_32_);
 assign n_209 = ~(R_15_15_ & T_14_32_);
 assign n_208 = ~(R_15_10_ & T_14_32_);
 assign n_207 = ~(R_15_13_ & T_14_32_);
 assign n_206 = ~(R_15_9_ & T_14_32_);
 assign n_205 = ~(R_15_1_ & T_14_32_);
 assign n_204 = ~(R_15_8_ & T_14_32_);
 assign n_203 = ~(R_15_12_ & T_14_32_);
 assign n_202 = ~(R_15_7_ & T_14_32_);
 assign n_201 = ~(R_15_6_ & T_14_32_);
 assign n_200 = ~(R_15_11_ & T_14_32_);
 assign n_199 = ~(R_15_5_ & T_14_32_);
 assign n_198 = (R_15_14_ & T_14_32_);
 assign R_14_16_ = ~(n_209 & (~T_14_16_ | T_14_32_));
 assign n_197 = ~(T_14_32_ & R_15_16_);
 assign n_196 = ~(T_14_32_ & n_1187);
 assign R_14_0_ = ~(n_196 & (~n_1191 | T_14_32_));
 assign n_195 = ~(T_14_32_ & R_15_2_);
 assign R_14_10_ = ~(n_206 & (~T_14_10_ | T_14_32_));
 assign R_14_14_ = ~(n_207 & (~T_14_14_ | T_14_32_));
 assign R_14_3_ = ~(n_195 & (~T_14_3_ | T_14_32_));
 assign R_14_2_ = ~(n_205 & (~T_14_2_ | T_14_32_));
 assign R_14_7_ = ~(n_201 & (~T_14_7_ | T_14_32_));
 assign n_194 = ~(n_983 & ~n_976);
 assign R_14_13_ = ~(n_203 & (~T_14_13_ | T_14_32_));
 assign n_193 = ~(T_14_32_ & R_15_3_);
 assign R_14_11_ = ~(n_982 & (~n_974 | n_976));
 assign R_14_1_ = ~(n_192 & (~T_14_1_ | T_14_32_));
 assign n_192 = ~(T_14_32_ & R_15_0_);
 assign R_14_6_ = ~(n_199 & (~T_14_6_ | T_14_32_));
 assign R_14_5_ = ~(n_210 & (~T_14_5_ | T_14_32_));
 assign R_14_4_ = ~(n_193 & (~T_14_4_ | T_14_32_));
 assign R_14_12_ = ~(n_200 & (~T_14_12_ | T_14_32_));
 assign R_14_9_ = ~(n_204 & (~T_14_9_ | T_14_32_));
 assign R_14_8_ = ~(n_202 & (~T_14_8_ | T_14_32_));
 assign R_14_17_ = ~(n_981 & (~n_975 | n_976));
 assign R_15_13_ = ~(n_184 & ~(R_16_12_ & n_171));
 assign R_15_0_ = ~(n_170 & (~n_1119 | T_15_32_));
 assign R_15_14_ = ~(n_178 & n_179);
 assign R_15_8_ = ~(n_169 & n_183);
 assign n_191 = ~(R_16_0_ & T_15_32_);
 assign n_190 = ~(R_16_15_ & n_173);
 assign n_189 = ~(R_16_9_ & n_176);
 assign n_188 = ~(R_16_2_ & T_15_32_);
 assign n_187 = ~(R_16_3_ & T_15_32_);
 assign n_186 = ~(R_16_1_ & T_15_32_);
 assign n_185 = ~(R_16_8_ & n_176);
 assign n_184 = ~(n_174 & T_15_13_);
 assign n_183 = ~(R_16_7_ & n_176);
 assign n_182 = ~(R_16_11_ & n_176);
 assign n_181 = ~(R_16_6_ & T_15_32_);
 assign n_180 = ~(R_16_5_ & T_15_32_);
 assign n_179 = ~(R_16_13_ & n_171);
 assign n_178 = ~(n_174 & T_15_14_);
 assign n_177 = ~(R_16_4_ & T_15_32_);
 assign n_176 = ~n_175;
 assign n_175 = ~T_15_32_;
 assign n_173 = ~n_174;
 assign n_174 = ~T_15_32_;
 assign n_171 = ~n_172;
 assign n_172 = ~T_15_32_;
 assign n_170 = ~(T_15_32_ & n_1111);
 assign R_15_3_ = ~(n_188 & (~T_15_3_ | T_15_32_));
 assign R_15_6_ = ~(n_180 & (~T_15_6_ | T_15_32_));
 assign n_169 = ~(n_174 & T_15_8_);
 assign R_15_2_ = ~(n_186 & (~T_15_2_ | T_15_32_));
 assign R_15_10_ = ~(n_189 & (~T_15_10_ | n_176));
 assign n_168 = ~(n_173 & R_16_14_);
 assign R_15_7_ = ~(n_181 & (~T_15_7_ | T_15_32_));
 assign R_15_9_ = ~(n_185 & (~T_15_9_ | n_171));
 assign n_167 = ~(n_171 & R_16_10_);
 assign R_15_1_ = ~(n_191 & (~T_15_1_ | T_15_32_));
 assign R_15_15_ = ~(n_168 & (~T_15_15_ | n_173));
 assign R_15_12_ = ~(n_182 & (~T_15_12_ | n_176));
 assign R_15_16_ = ~(n_190 & (~T_15_16_ | n_173));
 assign R_15_5_ = ~(n_177 & (~T_15_5_ | T_15_32_));
 assign R_15_4_ = ~(n_187 & (~T_15_4_ | T_15_32_));
 assign R_15_11_ = ~(n_167 & (~T_15_11_ | n_173));
 assign R_16_8_ = ~(n_161 & (~T_16_8_ | T_16_32_));
 assign R_16_15_ = ~(n_159 & ~n_149);
 assign R_16_11_ = ~(n_157 & n_158);
 assign R_16_13_ = ~(n_154 & n_150);
 assign R_16_7_ = ~(n_160 & (~T_16_7_ | T_16_32_));
 assign R_16_5_ = ~(n_155 & (~T_16_5_ | T_16_32_));
 assign R_16_4_ = ~(n_152 & (~T_16_4_ | T_16_32_));
 assign n_166 = ~(R_17_13_ & T_16_32_);
 assign n_165 = ~(R_17_8_ & T_16_32_);
 assign n_164 = ~(R_17_1_ & T_16_32_);
 assign n_163 = ~(R_17_11_ & T_16_32_);
 assign n_162 = ~(R_17_0_ & T_16_32_);
 assign n_161 = ~(R_17_7_ & T_16_32_);
 assign n_160 = ~(R_17_6_ & T_16_32_);
 assign n_159 = ~(n_151 & T_16_15_);
 assign n_158 = ~(R_17_10_ & T_16_32_);
 assign n_157 = ~(n_151 & T_16_11_);
 assign n_156 = ~(R_17_5_ & T_16_32_);
 assign n_155 = ~(R_17_4_ & T_16_32_);
 assign n_154 = ~(n_151 & T_16_13_);
 assign n_153 = ~(R_17_9_ & T_16_32_);
 assign n_152 = ~(R_17_3_ & T_16_32_);
 assign n_151 = ~T_16_32_;
 assign n_150 = ~(T_16_32_ & R_17_12_);
 assign R_16_3_ = ~(n_147 & (~T_16_3_ | T_16_32_));
 assign n_149 = ~(n_151 | ~R_17_14_);
 assign R_16_9_ = ~(n_165 & (~T_16_9_ | T_16_32_));
 assign R_16_2_ = ~(n_164 & (~T_16_2_ | T_16_32_));
 assign R_16_1_ = ~(n_162 & (~T_16_1_ | T_16_32_));
 assign R_16_0_ = ~(n_148 & (~n_1106 | T_16_32_));
 assign R_16_14_ = ~(n_166 & (~T_16_14_ | T_16_32_));
 assign R_16_6_ = ~(n_156 & (~T_16_6_ | T_16_32_));
 assign R_16_10_ = ~(n_153 & (~T_16_10_ | T_16_32_));
 assign R_16_12_ = ~(n_163 & (~T_16_12_ | T_16_32_));
 assign n_148 = ~(T_16_32_ & n_1084);
 assign n_147 = ~(T_16_32_ & R_17_2_);
 assign R_17_10_ = ~(n_137 & (~T_17_10_ | T_17_32_));
 assign R_17_11_ = ~(n_146 & ~(R_18_10_ & T_17_32_));
 assign R_17_8_ = ~(n_127 & n_144);
 assign R_17_7_ = ~(n_142 & (~T_17_7_ | T_17_32_));
 assign R_17_14_ = ~(n_138 & ~n_145);
 assign R_17_9_ = ~(n_133 & (T_17_32_ | n_131));
 assign R_17_5_ = ~(n_136 & (~T_17_5_ | T_17_32_));
 assign R_17_13_ = ~(n_132 & ~n_129);
 assign R_17_6_ = ~(n_139 & (~T_17_6_ | T_17_32_));
 assign R_17_4_ = ~(n_135 & (~T_17_4_ | T_17_32_));
 assign R_17_3_ = ~(n_140 & (~T_17_3_ | T_17_32_));
 assign R_17_2_ = ~(n_141 & (~T_17_2_ | T_17_32_));
 assign n_146 = ~(n_130 & T_17_11_);
 assign n_145 = ~(n_130 | ~R_18_13_);
 assign n_144 = ~(R_18_7_ & T_17_32_);
 assign n_143 = ~(R_18_0_ & T_17_32_);
 assign n_142 = ~(R_18_6_ & T_17_32_);
 assign n_141 = ~(R_18_1_ & T_17_32_);
 assign n_140 = ~(R_18_2_ & T_17_32_);
 assign n_139 = ~(R_18_5_ & T_17_32_);
 assign n_138 = ~(T_17_14_ & ~T_17_32_);
 assign n_137 = ~(R_18_9_ & T_17_32_);
 assign n_136 = ~(R_18_4_ & T_17_32_);
 assign n_135 = ~(R_18_3_ & T_17_32_);
 assign n_134 = ~(R_18_11_ & T_17_32_);
 assign n_133 = ~(R_18_8_ & T_17_32_);
 assign n_132 = ~(T_17_13_ & ~T_17_32_);
 assign n_131 = ~T_17_9_;
 assign n_130 = ~T_17_32_;
 assign n_129 = (R_18_12_ & T_17_32_);
 assign R_17_12_ = ~(n_134 & (~T_17_12_ | T_17_32_));
 assign n_128 = ~(T_17_32_ & n_1056);
 assign n_127 = ~(n_130 & T_17_8_);
 assign R_17_1_ = ~(n_143 & (~T_17_1_ | T_17_32_));
 assign R_17_0_ = ~(n_128 & (~T_17_0_ | T_17_32_));
 assign R_18_5_ = ~(n_117 & (~T_18_5_ | T_18_32_));
 assign R_18_6_ = ~(n_122 & (~T_18_6_ | T_18_32_));
 assign R_18_13_ = ~(n_120 & ~n_113);
 assign R_18_12_ = ~(n_125 & (T_18_32_ | n_114));
 assign R_18_11_ = ~(n_111 & ~(n_994 & T_18_32_));
 assign R_18_3_ = ~(n_121 & (~T_18_3_ | T_18_32_));
 assign R_18_4_ = ~(n_118 & (~T_18_4_ | T_18_32_));
 assign n_126 = ~(n_996 & T_18_32_);
 assign n_125 = ~(n_992 & T_18_32_);
 assign n_124 = ~(n_1013 & T_18_32_);
 assign n_123 = ~(n_1016 & T_18_32_);
 assign n_122 = ~(n_989 & T_18_32_);
 assign n_121 = ~(n_1003 & T_18_32_);
 assign n_120 = ~(T_18_13_ & ~T_18_32_);
 assign n_119 = ~(n_1008 & T_18_32_);
 assign n_118 = ~(n_1004 & T_18_32_);
 assign n_117 = ~(n_987 & T_18_32_);
 assign n_116 = ~(n_999 & T_18_32_);
 assign n_115 = ~(n_1000 & T_18_32_);
 assign n_114 = ~T_18_12_;
 assign n_113 = (n_995 & T_18_32_);
 assign R_18_0_ = ~(n_112 & (~n_1134 | T_18_32_));
 assign R_18_8_ = ~(n_116 & (~T_18_8_ | T_18_32_));
 assign R_18_2_ = ~(n_115 & (~T_18_2_ | T_18_32_));
 assign n_112 = ~(T_18_32_ & n_1121);
 assign R_18_10_ = ~(n_123 & (~T_18_10_ | T_18_32_));
 assign n_111 = ~(T_18_11_ & ~T_18_32_);
 assign R_18_7_ = ~(n_124 & (~T_18_7_ | T_18_32_));
 assign R_18_9_ = ~(n_126 & (~T_18_9_ | T_18_32_));
 assign R_18_1_ = ~(n_119 & (~T_18_1_ | T_18_32_));
 assign R_19_12_ = ~(n_102 & ~n_105);
 assign R_19_9_ = ~(n_100 & ~n_108);
 assign R_19_5_ = ~(n_107 & (~T_19_5_ | T_19_32_));
 assign R_19_0_ = ~(n_95 & (~T_19_0_ | T_19_32_));
 assign n_110 = ~(R_20_10_ & T_19_32_);
 assign n_109 = ~(R_20_5_ & T_19_32_);
 assign n_108 = ~(n_96 | ~R_20_8_);
 assign n_107 = ~(R_20_4_ & T_19_32_);
 assign n_106 = ~(R_20_7_ & T_19_32_);
 assign n_105 = ~(n_96 | ~R_20_11_);
 assign n_104 = ~(R_20_1_ & T_19_32_);
 assign n_103 = ~(R_20_3_ & T_19_32_);
 assign n_102 = ~(n_96 & T_19_12_);
 assign n_101 = ~(R_20_2_ & T_19_32_);
 assign n_100 = ~(n_96 & T_19_9_);
 assign n_99 = ~(R_20_9_ & T_19_32_);
 assign n_98 = ~(R_20_6_ & T_19_32_);
 assign n_97 = ~(R_20_0_ & T_19_32_);
 assign n_96 = ~T_19_32_;
 assign R_19_2_ = ~(n_104 & (~T_19_2_ | T_19_32_));
 assign R_19_4_ = ~(n_103 & (~T_19_4_ | T_19_32_));
 assign n_95 = ~(T_19_32_ & n_1024);
 assign R_19_11_ = ~(n_110 & (~T_19_11_ | T_19_32_));
 assign R_19_3_ = ~(n_101 & (~T_19_3_ | T_19_32_));
 assign R_19_1_ = ~(n_97 & (~T_19_1_ | T_19_32_));
 assign R_19_10_ = ~(n_99 & (~T_19_10_ | T_19_32_));
 assign R_19_8_ = ~(n_106 & (~T_19_8_ | T_19_32_));
 assign R_19_7_ = ~(n_98 & (~T_19_7_ | T_19_32_));
 assign R_19_6_ = ~(n_109 & (~T_19_6_ | T_19_32_));
 assign R_20_11_ = ~(n_81 & ~n_83);
 assign R_20_5_ = ~(n_93 & (~T_20_5_ | T_20_32_));
 assign R_20_4_ = ~(n_90 & (~T_20_4_ | T_20_32_));
 assign R_20_7_ = ~(n_92 & (~T_20_7_ | T_20_32_));
 assign R_20_3_ = ~(n_85 & (~T_20_3_ | T_20_32_));
 assign R_20_2_ = ~(n_89 & (~T_20_2_ | T_20_32_));
 assign R_20_9_ = ~(n_87 & (T_20_32_ | n_84));
 assign R_20_6_ = ~(n_86 & (~T_20_6_ | T_20_32_));
 assign R_20_0_ = ~(n_82 & (~T_20_0_ | T_20_32_));
 assign n_94 = ~(R_21_9_ & T_20_32_);
 assign n_93 = ~(R_21_4_ & T_20_32_);
 assign n_92 = ~(R_21_6_ & T_20_32_);
 assign n_91 = ~(R_21_7_ & T_20_32_);
 assign n_90 = ~(R_21_3_ & T_20_32_);
 assign n_89 = ~(R_21_1_ & T_20_32_);
 assign n_88 = ~(R_21_0_ & T_20_32_);
 assign n_87 = ~(R_21_8_ & T_20_32_);
 assign n_86 = ~(R_21_5_ & T_20_32_);
 assign n_85 = ~(R_21_2_ & T_20_32_);
 assign n_84 = ~T_20_9_;
 assign n_83 = (R_21_10_ & T_20_32_);
 assign R_20_8_ = ~(n_91 & (~T_20_8_ | T_20_32_));
 assign n_82 = ~(T_20_32_ & n_1109);
 assign R_20_10_ = ~(n_94 & (~T_20_10_ | T_20_32_));
 assign R_20_1_ = ~(n_88 & (~T_20_1_ | T_20_32_));
 assign n_81 = ~(T_20_11_ & ~T_20_32_);
 assign R_21_4_ = ~(n_79 & (~T_21_4_ | T_21_32_));
 assign R_21_7_ = ~(n_75 & ~(R_22_6_ & T_21_32_));
 assign R_21_10_ = ~(n_73 & ~n_65);
 assign R_21_3_ = ~(n_77 & (~T_21_3_ | T_21_32_));
 assign R_21_6_ = ~(n_80 & (T_21_32_ | n_70));
 assign R_21_2_ = ~(n_78 & (~T_21_2_ | T_21_32_));
 assign R_21_1_ = ~(n_72 & (~T_21_1_ | T_21_32_));
 assign R_21_9_ = ~(n_74 & ~n_67);
 assign R_21_8_ = ~(n_71 & (T_21_32_ | n_69));
 assign R_21_5_ = ~(n_76 & (~T_21_5_ | T_21_32_));
 assign R_21_0_ = ~(n_66 & (~T_21_0_ | T_21_32_));
 assign n_80 = ~(R_22_5_ & T_21_32_);
 assign n_79 = ~(R_22_3_ & T_21_32_);
 assign n_78 = ~(R_22_1_ & T_21_32_);
 assign n_77 = ~(R_22_2_ & T_21_32_);
 assign n_76 = ~(R_22_4_ & T_21_32_);
 assign n_75 = ~(n_68 & T_21_7_);
 assign n_74 = ~(n_68 & T_21_9_);
 assign n_73 = ~(n_68 & T_21_10_);
 assign n_72 = ~(R_22_0_ & T_21_32_);
 assign n_71 = ~(R_22_7_ & T_21_32_);
 assign n_70 = ~T_21_6_;
 assign n_69 = ~T_21_8_;
 assign n_68 = ~T_21_32_;
 assign n_67 = (R_22_8_ & T_21_32_);
 assign n_66 = ~(T_21_32_ & n_1018);
 assign n_65 = ~(n_68 | ~R_22_9_);
 assign R_22_3_ = ~(n_61 & (~T_22_3_ | T_22_32_));
 assign R_22_6_ = ~(n_60 & (~T_22_6_ | T_22_32_));
 assign R_22_9_ = ~(n_52 & ~n_54);
 assign R_22_2_ = ~(n_59 & (~T_22_2_ | T_22_32_));
 assign R_22_5_ = ~(n_64 & (~T_22_5_ | T_22_32_));
 assign R_22_8_ = ~(n_62 & (T_22_32_ | n_55));
 assign R_22_1_ = ~(n_63 & (~T_22_1_ | T_22_32_));
 assign R_22_7_ = ~(n_58 & (T_22_32_ | n_56));
 assign R_22_4_ = ~(n_57 & (~T_22_4_ | T_22_32_));
 assign n_64 = ~(R_23_4_ & T_22_32_);
 assign n_63 = ~(R_23_0_ & T_22_32_);
 assign n_62 = ~(R_23_7_ & T_22_32_);
 assign n_61 = ~(R_23_2_ & T_22_32_);
 assign n_60 = ~(R_23_5_ & T_22_32_);
 assign n_59 = ~(R_23_1_ & T_22_32_);
 assign n_58 = ~(R_23_6_ & T_22_32_);
 assign n_57 = ~(R_23_3_ & T_22_32_);
 assign n_56 = ~T_22_7_;
 assign n_55 = ~T_22_8_;
 assign n_54 = (R_23_8_ & T_22_32_);
 assign n_53 = ~(T_22_32_ & n_1057);
 assign R_22_0_ = ~(n_53 & (~T_22_0_ | T_22_32_));
 assign n_52 = ~(T_22_9_ & ~T_22_32_);
 assign R_23_5_ = ~(n_48 & (~T_23_5_ | T_23_32_));
 assign R_23_8_ = ~(n_50 & (~T_23_8_ | T_23_32_));
 assign R_23_0_ = ~(n_46 & n_40);
 assign n_51 = ~(R_24_6_ & T_23_32_);
 assign n_50 = ~(R_24_7_ & T_23_32_);
 assign n_49 = ~(R_24_1_ & T_23_32_);
 assign n_48 = ~(R_24_4_ & T_23_32_);
 assign n_47 = ~(R_24_3_ & T_23_32_);
 assign n_46 = ~(n_41 & ~n_1022);
 assign n_45 = ~(R_24_0_ & T_23_32_);
 assign n_44 = ~(R_24_5_ & T_23_32_);
 assign n_43 = ~(R_24_2_ & T_23_32_);
 assign n_42 = ~T_23_0_;
 assign n_41 = ~T_23_32_;
 assign R_23_1_ = ~(n_45 & (~T_23_1_ | T_23_32_));
 assign n_40 = ~(T_23_32_ & n_1017);
 assign R_23_2_ = ~(n_49 & (~T_23_2_ | T_23_32_));
 assign R_23_7_ = ~(n_51 & (~T_23_7_ | T_23_32_));
 assign R_23_6_ = ~(n_44 & (~T_23_6_ | T_23_32_));
 assign R_23_4_ = ~(n_47 & (~T_23_4_ | T_23_32_));
 assign R_23_3_ = ~(n_43 & (~T_23_3_ | T_23_32_));
 assign R_24_1_ = ~(n_1233 & (~n_1081 | n_1021));
 assign R_24_4_ = ~(n_1023 & n_1107);
 assign R_24_5_ = ~(n_1108 & (n_1021 | n_1078));
 assign R_24_6_ = ~(n_1079 & (n_1021 | n_32));
 assign R_24_3_ = ~(n_1043 & (~n_1290 | n_1021));
 assign R_24_2_ = ~(n_1082 & (~n_1020 | n_1021));
 assign n_39 = ~(R_25_0_ & T_24_32_);
 assign n_38 = ~(R_25_5_ & T_24_32_);
 assign n_37 = ~(R_25_6_ & T_24_32_);
 assign n_36 = ~(R_25_3_ & T_24_32_);
 assign n_35 = ~(R_25_2_ & T_24_32_);
 assign n_34 = ~(R_25_4_ & T_24_32_);
 assign n_33 = ~(R_25_1_ & T_24_32_);
 assign n_32 = ~n_1054;
 assign n_31 = ~T_24_5_;
 assign n_30 = ~(T_24_32_ & {in2[24]});
 assign R_24_0_ = ~(n_1053 & (~n_1207 | n_1021));
 assign R_24_7_ = ~(n_1117 & (~n_1080 | n_1021));
 assign n_29 = ~(T_24_4_ & ~T_24_32_);
 assign n_28 = ~(R_26_5_ & T_25_32_);
 assign n_27 = ~(R_26_4_ & T_25_32_);
 assign n_26 = ~(R_26_3_ & T_25_32_);
 assign n_25 = ~(R_26_1_ & T_25_32_);
 assign n_24 = ~(R_26_2_ & T_25_32_);
 assign n_23 = ~(R_26_0_ & T_25_32_);
 assign n_22 = ~(T_25_32_ & {in2[25]});
 assign R_25_0_ = ~(n_22 & (~T_25_0_ | T_25_32_));
 assign R_25_3_ = ~(n_24 & (~T_25_3_ | T_25_32_));
 assign R_25_4_ = ~(n_26 & (~T_25_4_ | T_25_32_));
 assign R_25_6_ = ~(n_28 & (~T_25_6_ | T_25_32_));
 assign R_25_1_ = ~(n_23 & (~T_25_1_ | T_25_32_));
 assign R_25_2_ = ~(n_25 & (~T_25_2_ | T_25_32_));
 assign R_25_5_ = ~(n_27 & (~T_25_5_ | T_25_32_));
 assign R_26_1_ = ~(n_19 & (~T_26_1_ | T_26_32_));
 assign R_26_3_ = ~(n_18 & (~T_26_3_ | T_26_32_));
 assign n_21 = ~(R_27_3_ & T_26_32_);
 assign n_20 = ~(R_27_1_ & T_26_32_);
 assign n_19 = ~(R_27_0_ & T_26_32_);
 assign n_18 = ~(R_27_2_ & T_26_32_);
 assign n_17 = ~(T_26_32_ & {in2[26]});
 assign R_26_5_ = ((T_26_5_ & ~T_26_32_) | (R_27_4_ & T_26_32_));
 assign R_26_2_ = ~(n_20 & (~T_26_2_ | T_26_32_));
 assign R_26_0_ = ~(n_17 & (~T_26_0_ | T_26_32_));
 assign R_26_4_ = ~(n_21 & (~T_26_4_ | T_26_32_));
 assign R_27_4_ = ~(n_16 & (T_27_32_ | n_12));
 assign n_16 = ~(R_28_3_ & T_27_32_);
 assign n_15 = ~(R_28_2_ & T_27_32_);
 assign n_14 = ~(R_28_0_ & T_27_32_);
 assign n_13 = ~(R_28_1_ & T_27_32_);
 assign n_12 = ~T_27_4_;
 assign n_11 = ~(T_27_32_ & {in2[27]});
 assign R_27_3_ = ~(n_15 & (~T_27_3_ | T_27_32_));
 assign R_27_0_ = ~(n_11 & (~T_27_0_ | T_27_32_));
 assign R_27_1_ = ~(n_14 & (~T_27_1_ | T_27_32_));
 assign R_27_2_ = ~(n_13 & (~T_27_2_ | T_27_32_));
 assign n_10 = ~(R_29_2_ & T_28_32_);
 assign n_9 = ~(R_29_1_ & T_28_32_);
 assign n_8 = ~(R_29_0_ & T_28_32_);
 assign n_7 = ~(T_28_32_ & {in2[28]});
 assign R_28_2_ = ~(n_9 & (~T_28_2_ | T_28_32_));
 assign R_28_0_ = ~(n_7 & (~T_28_0_ | T_28_32_));
 assign R_28_1_ = ~(n_8 & (~T_28_1_ | T_28_32_));
 assign R_28_3_ = ~(n_10 & (~T_28_3_ | T_28_32_));
 assign R_29_2_ = ~(n_3 & n_6);
 assign n_6 = ~(R_30_1_ & T_29_32_);
 assign n_5 = ~(R_30_0_ & T_29_32_);
 assign R_29_1_ = ~(n_5 & (~T_29_1_ | T_29_32_));
 assign n_4 = ~(T_29_32_ & {in2[29]});
 assign R_29_0_ = ~(n_4 & (~T_29_0_ | T_29_32_));
 assign n_3 = ~(T_29_2_ & ~T_29_32_);
 assign R_30_1_ = ~(n_2 & (~T_30_1_ | T_30_32_));
 assign n_2 = ~(R_31_0_ & T_30_32_);
 assign n_1 = ~(T_30_32_ & {in2[30]});
 assign R_30_0_ = ~(n_1 & (~T_30_0_ | T_30_32_));
 assign n_0 = ~(T_31_32_ & {in2[31]});
 assign R_31_0_ = ~(n_0 & (~T_31_0_ | T_31_32_));
 assign T_31_32_ = ~(sub_230_64_n_27 & (sub_230_64_n_23 & sub_230_64_n_25));
 assign sub_230_64_n_27 = ~(sub_230_64_n_26 | (sub_230_64_n_18 | ~sub_230_64_n_4));
 assign sub_230_64_n_26 = ~(sub_230_64_n_0 & ~{in1[1]});
 assign sub_230_64_n_25 = ~(sub_230_64_n_24 | sub_230_64_n_22);
 assign sub_230_64_n_24 = ~(sub_230_64_n_3 & (sub_230_64_n_6 & (sub_230_64_n_10 & sub_230_64_n_17)));
 assign sub_230_64_n_23 = ~(sub_230_64_n_19 | sub_230_64_n_20);
 assign sub_230_64_n_22 = ~(sub_230_64_n_9 & (sub_230_64_n_7 & (sub_230_64_n_13 & sub_230_64_n_11)));
 assign T_31_0_ = ~(sub_230_64_n_16 & sub_230_64_n_0);
 assign sub_230_64_n_20 = ~(sub_230_64_n_14 & sub_230_64_n_15);
 assign sub_230_64_n_19 = ~(sub_230_64_n_2 & sub_230_64_n_12);
 assign sub_230_64_n_18 = ~(sub_230_64_n_5 & sub_230_64_n_8);
 assign sub_230_64_n_17 = ~({in1[14]} | {in1[15]});
 assign sub_230_64_n_16 = ~({in2[31]} & ~{in1[0]});
 assign sub_230_64_n_15 = ~({in1[28]} | {in1[29]});
 assign sub_230_64_n_14 = ~({in1[26]} | {in1[27]});
 assign sub_230_64_n_13 = ~({in1[10]} | {in1[11]});
 assign sub_230_64_n_12 = ~({in1[24]} | {in1[25]});
 assign sub_230_64_n_11 = ~({in1[12]} | {in1[13]});
 assign sub_230_64_n_10 = ~({in1[4]} | {in1[5]});
 assign sub_230_64_n_9 = ~({in1[8]} | {in1[9]});
 assign sub_230_64_n_8 = ~({in1[20]} | {in1[21]});
 assign sub_230_64_n_7 = ~({in1[30]} | {in1[31]});
 assign sub_230_64_n_6 = ~({in1[6]} | {in1[7]});
 assign sub_230_64_n_5 = ~({in1[18]} | {in1[19]});
 assign sub_230_64_n_4 = ~({in1[16]} | {in1[17]});
 assign sub_230_64_n_3 = ~({in1[2]} | {in1[3]});
 assign sub_230_64_n_2 = ~({in1[22]} | {in1[23]});
 assign sub_230_64_n_0 = ~({in1[0]} & ~{in2[31]});
 assign T_30_1_ = ~((sub_260_63_n_36 | R_31_0_) & ~(sub_260_63_n_36 & R_31_0_));
 assign sub_260_63_n_37 = ~(sub_260_63_n_32 | (sub_260_63_n_33 | sub_260_63_n_34));
 assign sub_260_63_n_36 = ~(sub_260_63_n_1 & sub_260_63_n_35);
 assign sub_260_63_n_35 = ~(sub_260_63_n_0 & ~{in1[1]});
 assign sub_260_63_n_34 = ~(sub_260_63_n_0 | ~{in1[1]});
 assign sub_260_63_n_33 = ~(sub_260_63_n_30 & sub_260_63_n_28);
 assign sub_260_63_n_32 = ~(sub_260_63_n_29 & sub_260_63_n_31);
 assign sub_260_63_n_31 = ~(sub_260_63_n_23 | sub_260_63_n_24);
 assign sub_260_63_n_30 = ~(sub_260_63_n_26 | sub_260_63_n_22);
 assign sub_260_63_n_29 = ~(sub_260_63_n_20 | sub_260_63_n_21);
 assign sub_260_63_n_28 = ~(sub_260_63_n_25 | ~sub_260_63_n_5);
 assign T_30_0_ = ~(sub_260_63_n_14 & sub_260_63_n_0);
 assign sub_260_63_n_26 = ~(sub_260_63_n_16 & sub_260_63_n_17);
 assign sub_260_63_n_25 = ~(sub_260_63_n_13 & sub_260_63_n_19);
 assign sub_260_63_n_24 = ~(sub_260_63_n_6 & sub_260_63_n_12);
 assign sub_260_63_n_23 = ~(sub_260_63_n_18 & sub_260_63_n_9);
 assign sub_260_63_n_22 = ~(sub_260_63_n_4 & sub_260_63_n_7);
 assign sub_260_63_n_21 = ~(sub_260_63_n_11 & sub_260_63_n_10);
 assign sub_260_63_n_20 = ~(sub_260_63_n_8 & sub_260_63_n_15);
 assign sub_260_63_n_19 = ~({in1[12]} | {in1[13]});
 assign sub_260_63_n_18 = ~({in1[22]} | {in1[23]});
 assign sub_260_63_n_17 = ~({in1[6]} | {in1[7]});
 assign sub_260_63_n_16 = ~({in1[4]} | {in1[5]});
 assign sub_260_63_n_15 = ~({in1[16]} | {in1[17]});
 assign sub_260_63_n_14 = ~({in2[30]} & ~{in1[0]});
 assign sub_260_63_n_13 = ~({in1[2]} | {in1[3]});
 assign sub_260_63_n_12 = ~({in1[28]} | {in1[29]});
 assign sub_260_63_n_11 = ~({in1[18]} | {in1[19]});
 assign sub_260_63_n_10 = ~({in1[20]} | {in1[21]});
 assign sub_260_63_n_9 = ~({in1[24]} | {in1[25]});
 assign sub_260_63_n_8 = ~({in1[10]} | {in1[11]});
 assign sub_260_63_n_7 = ~({in1[14]} | {in1[15]});
 assign sub_260_63_n_6 = ~({in1[26]} | {in1[27]});
 assign sub_260_63_n_5 = ~({in1[30]} | {in1[31]});
 assign sub_260_63_n_4 = ~({in1[8]} | {in1[9]});
 assign T_30_32_ = ~(sub_260_63_n_37 & (~sub_260_63_n_35 | R_31_0_));
 assign sub_260_63_n_1 = ~({in1[1]} & ~sub_260_63_n_0);
 assign sub_260_63_n_0 = ~({in1[0]} & ~{in2[30]});
 assign T_29_32_ = ~(sub_290_62_n_40 & (sub_290_62_n_1 | sub_290_62_n_37));
 assign T_29_2_ = ~((sub_290_62_n_39 | sub_290_62_n_5) & ~(sub_290_62_n_39 & sub_290_62_n_5));
 assign sub_290_62_n_40 = ~(sub_290_62_n_38 | sub_290_62_n_25);
 assign sub_290_62_n_39 = ~((sub_290_62_n_3 & sub_290_62_n_9) | ((sub_290_62_n_9 & sub_290_62_n_6) |
    (sub_290_62_n_6 & sub_290_62_n_3)));
 assign sub_290_62_n_38 = ~(sub_290_62_n_33 & (sub_290_62_n_34 & sub_290_62_n_36));
 assign sub_290_62_n_37 = ~(sub_290_62_n_35 | (~sub_290_62_n_6 & sub_290_62_n_8));
 assign sub_290_62_n_36 = ~(sub_290_62_n_30 | (sub_290_62_n_27 | sub_290_62_n_4));
 assign sub_290_62_n_35 = ~sub_290_62_n_3;
 assign sub_290_62_n_34 = ~(sub_290_62_n_28 | sub_290_62_n_29);
 assign sub_290_62_n_33 = ~(sub_290_62_n_31 | sub_290_62_n_26);
 assign T_29_0_ = ~(sub_290_62_n_17 & sub_290_62_n_3);
 assign sub_290_62_n_31 = ~(sub_290_62_n_19 & sub_290_62_n_20);
 assign sub_290_62_n_30 = ~(sub_290_62_n_18 & sub_290_62_n_11);
 assign sub_290_62_n_29 = ~(sub_290_62_n_15 & sub_290_62_n_12);
 assign sub_290_62_n_28 = ~(sub_290_62_n_16 & sub_290_62_n_13);
 assign sub_290_62_n_27 = ~(sub_290_62_n_22 & sub_290_62_n_10);
 assign sub_290_62_n_26 = ~(sub_290_62_n_23 & sub_290_62_n_21);
 assign sub_290_62_n_24 = ~({in1[13]} | {in1[14]});
 assign sub_290_62_n_23 = ~({in1[5]} | {in1[6]});
 assign sub_290_62_n_22 = ~({in1[21]} | {in1[22]});
 assign sub_290_62_n_21 = ~({in1[7]} | {in1[28]});
 assign sub_290_62_n_20 = ~({in1[25]} | {in1[26]});
 assign sub_290_62_n_19 = ~({in1[4]} | {in1[27]});
 assign sub_290_62_n_18 = ~({in1[17]} | {in1[18]});
 assign sub_290_62_n_17 = ~({in2[29]} & ~{in1[0]});
 assign sub_290_62_n_25 = ~(R_30_1_ | ~{in1[2]});
 assign sub_290_62_n_16 = ~({in1[8]} | {in1[31]});
 assign sub_290_62_n_15 = ~({in1[9]} | {in1[10]});
 assign sub_290_62_n_14 = ~({in1[3]} | {in1[16]});
 assign sub_290_62_n_13 = ~({in1[29]} | {in1[30]});
 assign sub_290_62_n_12 = ~({in1[11]} | {in1[12]});
 assign sub_290_62_n_11 = ~({in1[19]} | {in1[20]});
 assign sub_290_62_n_10 = ~({in1[23]} | {in1[24]});
 assign sub_290_62_n_9 = ~sub_290_62_n_8;
 assign sub_290_62_n_8 = ~R_30_0_;
 assign sub_290_62_n_6 = ~{in1[1]};
 assign sub_290_62_n_5 = ~(sub_290_62_n_25 | ~sub_290_62_n_2);
 assign sub_290_62_n_4 = ~(sub_290_62_n_14 & (sub_290_62_n_24 & ~{in1[15]}));
 assign sub_290_62_n_3 = ~({in1[0]} & ~{in2[29]});
 assign sub_290_62_n_2 = ~(R_30_1_ & ~{in1[2]});
 assign sub_290_62_n_1 = ~(sub_290_62_n_2 & (~sub_290_62_n_6 | sub_290_62_n_8));
 assign T_29_1_ = ~(sub_290_62_n_9 ^ ({in1[1]} ^ sub_290_62_n_3));
 assign T_28_32_ = ~(sub_320_61_n_39 & sub_320_61_n_45);
 assign T_28_3_ = ~((sub_320_61_n_44 | sub_320_61_n_4) & ~(sub_320_61_n_44 & sub_320_61_n_4));
 assign sub_320_61_n_45 = ~(sub_320_61_n_43 & ~sub_320_61_n_31);
 assign sub_320_61_n_44 = ~(sub_320_61_n_41 | ~sub_320_61_n_1);
 assign sub_320_61_n_43 = ~(sub_320_61_n_41 & ~sub_320_61_n_21);
 assign T_28_2_ = ~((sub_320_61_n_40 | sub_320_61_n_30) & ~(sub_320_61_n_40 & sub_320_61_n_30));
 assign sub_320_61_n_41 = ~(sub_320_61_n_38 | ~sub_320_61_n_0);
 assign sub_320_61_n_40 = ~sub_320_61_n_38;
 assign sub_320_61_n_39 = ~(sub_320_61_n_35 | sub_320_61_n_36);
 assign sub_320_61_n_38 = ~((sub_320_61_n_3 & R_29_0_) | ((R_29_0_ & sub_320_61_n_6) | (sub_320_61_n_6
    & sub_320_61_n_3)));
 assign T_28_1_ = ~(R_29_0_ ^ ({in1[1]} ^ sub_320_61_n_3));
 assign sub_320_61_n_36 = ~(sub_320_61_n_34 & ~sub_320_61_n_23);
 assign sub_320_61_n_35 = ~(sub_320_61_n_33 & sub_320_61_n_32);
 assign sub_320_61_n_34 = ~(sub_320_61_n_25 | sub_320_61_n_27);
 assign sub_320_61_n_33 = ~(sub_320_61_n_26 | sub_320_61_n_28);
 assign sub_320_61_n_32 = ~(sub_320_61_n_22 | sub_320_61_n_24);
 assign sub_320_61_n_31 = ~(sub_320_61_n_2 & (sub_320_61_n_1 | sub_320_61_n_21));
 assign sub_320_61_n_30 = ~(sub_320_61_n_1 & sub_320_61_n_0);
 assign T_28_0_ = ~(sub_320_61_n_3 & (~{in2[28]} | {in1[0]}));
 assign sub_320_61_n_28 = ~(sub_320_61_n_17 & sub_320_61_n_19);
 assign sub_320_61_n_27 = ~(sub_320_61_n_20 & sub_320_61_n_16);
 assign sub_320_61_n_26 = ~(sub_320_61_n_18 & sub_320_61_n_15);
 assign sub_320_61_n_25 = ~(sub_320_61_n_13 & sub_320_61_n_14);
 assign sub_320_61_n_24 = ~(sub_320_61_n_9 & sub_320_61_n_11);
 assign sub_320_61_n_23 = ~(sub_320_61_n_8 & sub_320_61_n_10);
 assign sub_320_61_n_22 = ~(sub_320_61_n_12 & sub_320_61_n_7);
 assign sub_320_61_n_20 = ~({in1[8]} | {in1[9]});
 assign sub_320_61_n_19 = ~({in1[18]} | {in1[19]});
 assign sub_320_61_n_18 = ~({in1[12]} | {in1[13]});
 assign sub_320_61_n_17 = ~({in1[16]} | {in1[17]});
 assign sub_320_61_n_16 = ~({in1[10]} | {in1[11]});
 assign sub_320_61_n_15 = ~({in1[14]} | {in1[15]});
 assign sub_320_61_n_21 = ~(R_29_2_ | ~{in1[3]});
 assign sub_320_61_n_14 = ~({in1[6]} | {in1[7]});
 assign sub_320_61_n_13 = ~({in1[4]} | {in1[5]});
 assign sub_320_61_n_12 = ~({in1[20]} | {in1[21]});
 assign sub_320_61_n_11 = ~({in1[26]} | {in1[27]});
 assign sub_320_61_n_10 = ~({in1[30]} | {in1[31]});
 assign sub_320_61_n_9 = ~({in1[24]} | {in1[25]});
 assign sub_320_61_n_8 = ~({in1[28]} | {in1[29]});
 assign sub_320_61_n_7 = ~({in1[22]} | {in1[23]});
 assign sub_320_61_n_6 = ~{in1[1]};
 assign sub_320_61_n_4 = ~(sub_320_61_n_21 | ~sub_320_61_n_2);
 assign sub_320_61_n_3 = ~({in1[0]} & ~{in2[28]});
 assign sub_320_61_n_2 = ~(R_29_2_ & ~{in1[3]});
 assign sub_320_61_n_1 = ~(R_29_1_ & ~{in1[2]});
 assign sub_320_61_n_0 = ~({in1[2]} & ~R_29_1_);
 assign T_27_32_ = ~(sub_350_60_n_47 & sub_350_60_n_56);
 assign T_27_4_ = ((sub_350_60_n_54 & sub_350_60_n_38) | ~(sub_350_60_n_54 | sub_350_60_n_38));
 assign T_27_3_ = ((sub_350_60_n_55 & sub_350_60_n_39) | ~(sub_350_60_n_55 | sub_350_60_n_39));
 assign sub_350_60_n_56 = ((sub_350_60_n_40 & sub_350_60_n_34) | ~(sub_350_60_n_51 | sub_350_60_n_43));
 assign sub_350_60_n_55 = ~(sub_350_60_n_52 | ~sub_350_60_n_0);
 assign sub_350_60_n_54 = ~(sub_350_60_n_41 | (sub_350_60_n_49 & sub_350_60_n_37));
 assign T_27_2_ = ~((sub_350_60_n_50 | sub_350_60_n_3) & ~(sub_350_60_n_50 & sub_350_60_n_3));
 assign sub_350_60_n_52 = ~sub_350_60_n_51;
 assign sub_350_60_n_51 = ~(sub_350_60_n_49 & ~sub_350_60_n_4);
 assign sub_350_60_n_50 = ~sub_350_60_n_49;
 assign sub_350_60_n_49 = ((sub_350_60_n_2 & R_28_0_) | ((R_28_0_ & sub_350_60_n_7) | (sub_350_60_n_7
    & sub_350_60_n_2)));
 assign T_27_1_ = (R_28_0_ ^ (sub_350_60_n_7 ^ sub_350_60_n_2));
 assign sub_350_60_n_47 = ~(sub_350_60_n_46 | sub_350_60_n_1);
 assign sub_350_60_n_46 = ~(sub_350_60_n_45 & (sub_350_60_n_42 & sub_350_60_n_44));
 assign sub_350_60_n_45 = ~(sub_350_60_n_30 | sub_350_60_n_31);
 assign sub_350_60_n_44 = ~(sub_350_60_n_32 | sub_350_60_n_29);
 assign sub_350_60_n_43 = ~(sub_350_60_n_34 & sub_350_60_n_27);
 assign sub_350_60_n_42 = ~(sub_350_60_n_33 | sub_350_60_n_28);
 assign sub_350_60_n_41 = ~(sub_350_60_n_19 & (sub_350_60_n_0 | sub_350_60_n_5));
 assign sub_350_60_n_40 = ~(sub_350_60_n_36 & (sub_350_60_n_0 | sub_350_60_n_5));
 assign sub_350_60_n_37 = ~(sub_350_60_n_4 | sub_350_60_n_5);
 assign sub_350_60_n_36 = ~(sub_350_60_n_18 | sub_350_60_n_20);
 assign T_27_0_ = ~(sub_350_60_n_15 & sub_350_60_n_2);
 assign sub_350_60_n_39 = ~(sub_350_60_n_18 | sub_350_60_n_5);
 assign sub_350_60_n_38 = ~(sub_350_60_n_20 | sub_350_60_n_1);
 assign sub_350_60_n_33 = ~(sub_350_60_n_22 & sub_350_60_n_13);
 assign sub_350_60_n_32 = ~(sub_350_60_n_12 & sub_350_60_n_11);
 assign sub_350_60_n_31 = ~(sub_350_60_n_17 & sub_350_60_n_25);
 assign sub_350_60_n_30 = ~(sub_350_60_n_21 & sub_350_60_n_26);
 assign sub_350_60_n_29 = ~(sub_350_60_n_23 & sub_350_60_n_24);
 assign sub_350_60_n_28 = ~(sub_350_60_n_16 & sub_350_60_n_14);
 assign sub_350_60_n_34 = ~({in1[6]} | ({in1[7]} | {in1[5]}));
 assign sub_350_60_n_27 = ~sub_350_60_n_5;
 assign sub_350_60_n_26 = ~({in1[10]} | {in1[11]});
 assign sub_350_60_n_25 = ~({in1[14]} | {in1[15]});
 assign sub_350_60_n_24 = ~({in1[30]} | {in1[31]});
 assign sub_350_60_n_23 = ~({in1[28]} | {in1[29]});
 assign sub_350_60_n_22 = ~({in1[16]} | {in1[17]});
 assign sub_350_60_n_21 = ~({in1[8]} | {in1[9]});
 assign sub_350_60_n_5 = ~(sub_350_60_n_10 | ~{in1[3]});
 assign sub_350_60_n_19 = ~sub_350_60_n_18;
 assign sub_350_60_n_17 = ~({in1[12]} | {in1[13]});
 assign sub_350_60_n_16 = ~({in1[20]} | {in1[21]});
 assign sub_350_60_n_15 = ~({in2[27]} & ~{in1[0]});
 assign sub_350_60_n_14 = ~({in1[22]} | {in1[23]});
 assign sub_350_60_n_13 = ~({in1[18]} | {in1[19]});
 assign sub_350_60_n_12 = ~({in1[24]} | {in1[25]});
 assign sub_350_60_n_11 = ~({in1[26]} | {in1[27]});
 assign sub_350_60_n_20 = ~({in1[4]} | sub_350_60_n_8);
 assign sub_350_60_n_18 = ~({in1[3]} | sub_350_60_n_9);
 assign sub_350_60_n_10 = ~sub_350_60_n_9;
 assign sub_350_60_n_9 = ~R_28_2_;
 assign sub_350_60_n_8 = ~R_28_3_;
 assign sub_350_60_n_7 = ~{in1[1]};
 assign sub_350_60_n_4 = ~(R_28_1_ | ~{in1[2]});
 assign sub_350_60_n_3 = ~(sub_350_60_n_4 | ~sub_350_60_n_0);
 assign sub_350_60_n_2 = ~({in1[0]} & ~{in2[27]});
 assign sub_350_60_n_1 = (sub_350_60_n_8 & {in1[4]});
 assign sub_350_60_n_0 = ~(R_28_1_ & ~{in1[2]});
 assign T_26_5_ = ((sub_380_59_n_61 & sub_380_59_n_41) | ~(sub_380_59_n_61 | sub_380_59_n_41));
 assign T_26_4_ = ((sub_380_59_n_63 & sub_380_59_n_42) | ~(sub_380_59_n_63 | sub_380_59_n_42));
 assign T_26_3_ = ~((sub_380_59_n_6 | sub_380_59_n_4) & ~(sub_380_59_n_6 & sub_380_59_n_4));
 assign T_26_32_ = ~(sub_380_59_n_55 & sub_380_59_n_62);
 assign sub_380_59_n_63 = ~(sub_380_59_n_48 | (sub_380_59_n_57 & sub_380_59_n_44));
 assign sub_380_59_n_62 = ~(sub_380_59_n_47 & (sub_380_59_n_45 & sub_380_59_n_59));
 assign sub_380_59_n_61 = ~(sub_380_59_n_52 & (sub_380_59_n_49 | sub_380_59_n_58));
 assign T_26_2_ = ~((sub_380_59_n_58 | sub_380_59_n_5) & ~(sub_380_59_n_58 & sub_380_59_n_5));
 assign sub_380_59_n_59 = ~(sub_380_59_n_57 & sub_380_59_n_44);
 assign sub_380_59_n_58 = ~sub_380_59_n_57;
 assign sub_380_59_n_57 = ((sub_380_59_n_3 & R_27_0_) | ((R_27_0_ & sub_380_59_n_11) | (sub_380_59_n_11
    & sub_380_59_n_3)));
 assign T_26_1_ = (R_27_0_ ^ (sub_380_59_n_11 ^ sub_380_59_n_3));
 assign sub_380_59_n_55 = ~(sub_380_59_n_54 | (sub_380_59_n_45 & sub_380_59_n_40));
 assign sub_380_59_n_54 = ~(sub_380_59_n_51 & (sub_380_59_n_50 & sub_380_59_n_53));
 assign sub_380_59_n_53 = ~(sub_380_59_n_46 | sub_380_59_n_32);
 assign sub_380_59_n_52 = ~(sub_380_59_n_22 | (sub_380_59_n_43 & sub_380_59_n_38));
 assign sub_380_59_n_51 = ~(sub_380_59_n_33 | sub_380_59_n_37);
 assign sub_380_59_n_50 = ~(sub_380_59_n_34 | sub_380_59_n_36);
 assign sub_380_59_n_49 = ~(sub_380_59_n_43 & ~sub_380_59_n_8);
 assign sub_380_59_n_48 = ~sub_380_59_n_47;
 assign sub_380_59_n_47 = ~(sub_380_59_n_38 & ~sub_380_59_n_20);
 assign sub_380_59_n_46 = ~(sub_380_59_n_14 & (sub_380_59_n_13 & sub_380_59_n_27));
 assign sub_380_59_n_45 = ~(sub_380_59_n_39 & sub_380_59_n_2);
 assign sub_380_59_n_40 = ~(sub_380_59_n_1 & sub_380_59_n_2);
 assign sub_380_59_n_39 = ~(sub_380_59_n_21 & sub_380_59_n_23);
 assign sub_380_59_n_44 = ~(sub_380_59_n_8 | sub_380_59_n_20);
 assign sub_380_59_n_43 = ~(sub_380_59_n_20 | sub_380_59_n_31);
 assign sub_380_59_n_42 = ~(sub_380_59_n_22 | sub_380_59_n_31);
 assign sub_380_59_n_41 = ~(sub_380_59_n_23 & sub_380_59_n_2);
 assign sub_380_59_n_37 = ~(sub_380_59_n_30 & sub_380_59_n_24);
 assign sub_380_59_n_36 = ~(sub_380_59_n_28 & sub_380_59_n_17);
 assign T_26_0_ = ~(sub_380_59_n_16 & sub_380_59_n_3);
 assign sub_380_59_n_34 = ~(sub_380_59_n_29 & sub_380_59_n_26);
 assign sub_380_59_n_33 = ~(sub_380_59_n_15 & sub_380_59_n_25);
 assign sub_380_59_n_32 = ~(sub_380_59_n_18 & sub_380_59_n_19);
 assign sub_380_59_n_38 = ~(sub_380_59_n_7 & sub_380_59_n_0);
 assign sub_380_59_n_30 = ~({in1[14]} | {in1[15]});
 assign sub_380_59_n_29 = ~({in1[18]} | {in1[19]});
 assign sub_380_59_n_28 = ~({in1[22]} | {in1[23]});
 assign sub_380_59_n_27 = ~({in1[30]} | {in1[31]});
 assign sub_380_59_n_26 = ~({in1[20]} | {in1[21]});
 assign sub_380_59_n_25 = ~({in1[12]} | {in1[13]});
 assign sub_380_59_n_24 = ~({in1[16]} | {in1[17]});
 assign sub_380_59_n_31 = ~(R_27_3_ | ~{in1[4]});
 assign sub_380_59_n_8 = ~(R_27_1_ | ~{in1[2]});
 assign sub_380_59_n_22 = ~sub_380_59_n_21;
 assign sub_380_59_n_19 = ~({in1[28]} | {in1[29]});
 assign sub_380_59_n_18 = ~({in1[26]} | {in1[27]});
 assign sub_380_59_n_17 = ~({in1[24]} | {in1[25]});
 assign sub_380_59_n_16 = ~({in2[26]} & ~{in1[0]});
 assign sub_380_59_n_15 = ~({in1[10]} | {in1[11]});
 assign sub_380_59_n_14 = ~({in1[6]} | {in1[7]});
 assign sub_380_59_n_13 = ~({in1[8]} | {in1[9]});
 assign sub_380_59_n_23 = ~(sub_380_59_n_10 & R_27_4_);
 assign sub_380_59_n_7 = ~(R_27_1_ & ~{in1[2]});
 assign sub_380_59_n_21 = ~(sub_380_59_n_12 & R_27_3_);
 assign sub_380_59_n_20 = ~(R_27_2_ | ~{in1[3]});
 assign sub_380_59_n_12 = ~{in1[4]};
 assign sub_380_59_n_11 = ~{in1[1]};
 assign sub_380_59_n_10 = ~{in1[5]};
 assign sub_380_59_n_6 = ~(sub_380_59_n_7 & (sub_380_59_n_8 | sub_380_59_n_58));
 assign sub_380_59_n_5 = ~(sub_380_59_n_8 | ~sub_380_59_n_7);
 assign sub_380_59_n_4 = ~(sub_380_59_n_0 & ~sub_380_59_n_20);
 assign sub_380_59_n_3 = ~({in1[0]} & ~{in2[26]});
 assign sub_380_59_n_2 = (R_27_4_ | sub_380_59_n_10);
 assign sub_380_59_n_1 = (R_27_3_ | sub_380_59_n_12);
 assign sub_380_59_n_0 = ~(R_27_2_ & ~{in1[3]});
 assign T_25_32_ = ~(sub_410_58_n_69 & sub_410_58_n_59);
 assign T_25_6_ = ((sub_410_58_n_12 & sub_410_58_n_6) | ~(sub_410_58_n_12 | sub_410_58_n_6));
 assign T_25_5_ = ((sub_410_58_n_9 & sub_410_58_n_7) | ~(sub_410_58_n_9 | sub_410_58_n_7));
 assign sub_410_58_n_69 = ~(sub_410_58_n_67 & ~sub_410_58_n_13);
 assign T_25_3_ = ~((sub_410_58_n_64 | sub_410_58_n_11) & ~(sub_410_58_n_64 & sub_410_58_n_11));
 assign sub_410_58_n_67 = ~(sub_410_58_n_65 & ~sub_410_58_n_48);
 assign T_25_4_ = ((sub_410_58_n_62 & sub_410_58_n_10) | ~(sub_410_58_n_62 | sub_410_58_n_10));
 assign sub_410_58_n_65 = ~(sub_410_58_n_60 | ~sub_410_58_n_49);
 assign sub_410_58_n_64 = ~(sub_410_58_n_25 | (~sub_410_58_n_35 & sub_410_58_n_5));
 assign T_25_2_ = ((sub_410_58_n_5 & sub_410_58_n_8) | ~(sub_410_58_n_5 | sub_410_58_n_8));
 assign sub_410_58_n_62 = ~sub_410_58_n_61;
 assign sub_410_58_n_61 = ~sub_410_58_n_60;
 assign sub_410_58_n_60 = ~(sub_410_58_n_51 | (sub_410_58_n_47 & (sub_410_58_n_4 & sub_410_58_n_57)));
 assign sub_410_58_n_59 = ~(sub_410_58_n_56 | ~sub_410_58_n_52);
 assign T_25_1_ = ((sub_410_58_n_46 & sub_410_58_n_55) | ~(sub_410_58_n_46 | sub_410_58_n_55));
 assign sub_410_58_n_57 = ~(sub_410_58_n_23 & sub_410_58_n_37);
 assign sub_410_58_n_56 = ~(sub_410_58_n_54 & sub_410_58_n_53);
 assign sub_410_58_n_55 = ~sub_410_58_n_23;
 assign sub_410_58_n_54 = ~(sub_410_58_n_44 | sub_410_58_n_42);
 assign sub_410_58_n_53 = ~(sub_410_58_n_45 | sub_410_58_n_39);
 assign sub_410_58_n_52 = ~(sub_410_58_n_40 | sub_410_58_n_41);
 assign sub_410_58_n_51 = ~(sub_410_58_n_2 & (sub_410_58_n_24 | sub_410_58_n_36));
 assign sub_410_58_n_50 = ~(sub_410_58_n_27 & (sub_410_58_n_38 | sub_410_58_n_34));
 assign sub_410_58_n_48 = ~sub_410_58_n_0;
 assign sub_410_58_n_49 = ~(sub_410_58_n_14 | sub_410_58_n_34);
 assign sub_410_58_n_47 = ~(sub_410_58_n_35 | sub_410_58_n_36);
 assign sub_410_58_n_45 = ~(sub_410_58_n_29 & sub_410_58_n_21);
 assign sub_410_58_n_44 = ~(sub_410_58_n_20 & sub_410_58_n_33);
 assign T_25_0_ = ~(sub_410_58_n_19 & sub_410_58_n_55);
 assign sub_410_58_n_42 = ~(sub_410_58_n_30 & sub_410_58_n_32);
 assign sub_410_58_n_41 = ~(sub_410_58_n_31 & sub_410_58_n_22);
 assign sub_410_58_n_40 = ~(sub_410_58_n_17 & sub_410_58_n_18);
 assign sub_410_58_n_39 = ~(sub_410_58_n_16 & sub_410_58_n_28);
 assign sub_410_58_n_46 = ~(sub_410_58_n_37 & sub_410_58_n_4);
 assign sub_410_58_n_33 = ~({in1[10]} | {in1[11]});
 assign sub_410_58_n_32 = ~({in1[14]} | {in1[15]});
 assign sub_410_58_n_31 = ~({in1[28]} | {in1[29]});
 assign sub_410_58_n_30 = ~({in1[12]} | {in1[13]});
 assign sub_410_58_n_29 = ~({in1[16]} | {in1[17]});
 assign sub_410_58_n_28 = ~({in1[22]} | {in1[23]});
 assign sub_410_58_n_38 = ~(R_26_3_ & ~{in1[4]});
 assign sub_410_58_n_37 = ~(R_26_0_ & ~{in1[1]});
 assign sub_410_58_n_36 = ~(R_26_2_ | ~{in1[3]});
 assign sub_410_58_n_14 = ~(R_26_3_ | ~{in1[4]});
 assign sub_410_58_n_35 = ~(R_26_1_ | ~{in1[2]});
 assign sub_410_58_n_34 = ~(R_26_4_ | ~{in1[5]});
 assign sub_410_58_n_25 = ~sub_410_58_n_24;
 assign sub_410_58_n_22 = ~({in1[30]} | {in1[31]});
 assign sub_410_58_n_21 = ~({in1[18]} | {in1[19]});
 assign sub_410_58_n_20 = ~({in1[8]} | {in1[9]});
 assign sub_410_58_n_19 = ~({in2[25]} & ~{in1[0]});
 assign sub_410_58_n_18 = ~({in1[26]} | {in1[27]});
 assign sub_410_58_n_17 = ~({in1[24]} | {in1[25]});
 assign sub_410_58_n_16 = ~({in1[20]} | {in1[21]});
 assign sub_410_58_n_27 = ~(R_26_4_ & ~{in1[5]});
 assign sub_410_58_n_26 = ~(R_26_5_ | ~{in1[6]});
 assign sub_410_58_n_24 = ~(R_26_1_ & ~{in1[2]});
 assign sub_410_58_n_23 = ~({in2[25]} | ~{in1[0]});
 assign sub_410_58_n_13 = (sub_410_58_n_1 | (sub_410_58_n_50 & sub_410_58_n_0));
 assign sub_410_58_n_12 = ~(sub_410_58_n_50 | (sub_410_58_n_49 & sub_410_58_n_61));
 assign sub_410_58_n_11 = ~(sub_410_58_n_36 | ~sub_410_58_n_2);
 assign sub_410_58_n_10 = ~(sub_410_58_n_14 | ~sub_410_58_n_38);
 assign sub_410_58_n_9 = ~(sub_410_58_n_38 & (sub_410_58_n_14 | sub_410_58_n_60));
 assign sub_410_58_n_8 = ~(sub_410_58_n_24 & ~sub_410_58_n_35);
 assign sub_410_58_n_7 = ~(sub_410_58_n_27 & ~sub_410_58_n_34);
 assign sub_410_58_n_6 = ~(sub_410_58_n_26 | ~sub_410_58_n_3);
 assign sub_410_58_n_5 = ~(sub_410_58_n_37 & (~sub_410_58_n_4 | sub_410_58_n_23));
 assign sub_410_58_n_4 = ~({in1[1]} & ~R_26_0_);
 assign sub_410_58_n_3 = ~(R_26_5_ & ~{in1[6]});
 assign sub_410_58_n_2 = ~(R_26_2_ & ~{in1[3]});
 assign sub_410_58_n_1 = ~(sub_410_58_n_3 | {in1[7]});
 assign sub_410_58_n_0 = ~(sub_410_58_n_26 | {in1[7]});
 assign T_24_7_ = ~((sub_440_57_n_80 | sub_440_57_n_9) & ~(sub_440_57_n_80 & sub_440_57_n_9));
 assign T_24_6_ = ~((sub_440_57_n_79 | sub_440_57_n_8) & ~(sub_440_57_n_79 & sub_440_57_n_8));
 assign T_24_5_ = ~((sub_440_57_n_78 | sub_440_57_n_49) & ~(sub_440_57_n_78 & sub_440_57_n_49));
 assign T_24_32_ = ~(sub_440_57_n_81 & sub_440_57_n_71);
 assign T_24_3_ = ((sub_440_57_n_76 & sub_440_57_n_52) | ~(sub_440_57_n_76 | sub_440_57_n_52));
 assign sub_440_57_n_81 = ~(sub_440_57_n_72 & (sub_440_57_n_63 & sub_440_57_n_73));
 assign sub_440_57_n_80 = ~(sub_440_57_n_66 | (~sub_440_57_n_57 & sub_440_57_n_74));
 assign sub_440_57_n_79 = ~(sub_440_57_n_59 | (~sub_440_57_n_46 & sub_440_57_n_74));
 assign sub_440_57_n_78 = ~(sub_440_57_n_25 | (~sub_440_57_n_24 & sub_440_57_n_74));
 assign T_24_4_ = ((sub_440_57_n_74 & sub_440_57_n_6) | ~(sub_440_57_n_74 | sub_440_57_n_6));
 assign sub_440_57_n_76 = ~(sub_440_57_n_34 & (~sub_440_57_n_27 | sub_440_57_n_69));
 assign T_24_2_ = ~((sub_440_57_n_70 | sub_440_57_n_53) & ~(sub_440_57_n_70 & sub_440_57_n_53));
 assign sub_440_57_n_74 = ~(sub_440_57_n_68 & ~sub_440_57_n_56);
 assign sub_440_57_n_73 = ~(sub_440_57_n_48 & (sub_440_57_n_12 | (sub_440_57_n_56 & sub_440_57_n_45)));
 assign sub_440_57_n_72 = ~(sub_440_57_n_67 & sub_440_57_n_60);
 assign sub_440_57_n_71 = (sub_440_57_n_39 & (sub_440_57_n_40 & sub_440_57_n_62));
 assign sub_440_57_n_70 = ~sub_440_57_n_69;
 assign sub_440_57_n_69 = ~(sub_440_57_n_7 | ~sub_440_57_n_26);
 assign sub_440_57_n_68 = ~sub_440_57_n_67;
 assign sub_440_57_n_67 = ~(sub_440_57_n_54 | ~sub_440_57_n_64);
 assign sub_440_57_n_66 = ~(sub_440_57_n_36 & (~sub_440_57_n_3 | sub_440_57_n_58));
 assign T_24_1_ = ~((sub_440_57_n_50 | sub_440_57_n_61) & ~(sub_440_57_n_50 & sub_440_57_n_61));
 assign sub_440_57_n_64 = ~(sub_440_57_n_21 & sub_440_57_n_26);
 assign sub_440_57_n_63 = ~(sub_440_57_n_55 | (sub_440_57_n_51 & sub_440_57_n_48));
 assign sub_440_57_n_62 = ~(sub_440_57_n_43 | (sub_440_57_n_44 | (sub_440_57_n_41 | sub_440_57_n_38)));
 assign sub_440_57_n_61 = ~sub_440_57_n_21;
 assign sub_440_57_n_60 = ~(sub_440_57_n_46 | sub_440_57_n_47);
 assign sub_440_57_n_59 = ~sub_440_57_n_58;
 assign sub_440_57_n_58 = ~(sub_440_57_n_51 | ~sub_440_57_n_11);
 assign sub_440_57_n_57 = ~(sub_440_57_n_45 & ~sub_440_57_n_22);
 assign sub_440_57_n_56 = ~(sub_440_57_n_0 & (sub_440_57_n_34 | sub_440_57_n_32));
 assign sub_440_57_n_55 = ~(sub_440_57_n_37 & (sub_440_57_n_36 | sub_440_57_n_23));
 assign sub_440_57_n_54 = ~(sub_440_57_n_27 & (sub_440_57_n_33 & sub_440_57_n_4));
 assign sub_440_57_n_53 = ~(sub_440_57_n_34 & sub_440_57_n_27);
 assign sub_440_57_n_52 = ~(sub_440_57_n_0 & sub_440_57_n_33);
 assign sub_440_57_n_51 = ~(sub_440_57_n_2 | sub_440_57_n_35);
 assign sub_440_57_n_50 = ~(sub_440_57_n_26 & sub_440_57_n_4);
 assign sub_440_57_n_49 = ~(sub_440_57_n_12 | sub_440_57_n_35);
 assign sub_440_57_n_47 = ~(sub_440_57_n_3 & sub_440_57_n_5);
 assign sub_440_57_n_48 = ~(sub_440_57_n_22 | sub_440_57_n_23);
 assign sub_440_57_n_44 = ~(sub_440_57_n_28 & sub_440_57_n_29);
 assign sub_440_57_n_43 = ~(sub_440_57_n_19 & sub_440_57_n_31);
 assign T_24_0_ = ~(sub_440_57_n_61 & (~{in2[24]} | {in1[0]}));
 assign sub_440_57_n_41 = ~(sub_440_57_n_18 & sub_440_57_n_30);
 assign sub_440_57_n_40 = ~({in1[28]} | ({in1[29]} | ({in1[30]} | {in1[31]})));
 assign sub_440_57_n_39 = ~({in1[24]} | ({in1[25]} | ({in1[26]} | {in1[27]})));
 assign sub_440_57_n_38 = ~(sub_440_57_n_20 & sub_440_57_n_17);
 assign sub_440_57_n_46 = ~(sub_440_57_n_10 & sub_440_57_n_1);
 assign sub_440_57_n_45 = ~(sub_440_57_n_24 | sub_440_57_n_35);
 assign sub_440_57_n_12 = ~sub_440_57_n_11;
 assign sub_440_57_n_33 = ~sub_440_57_n_32;
 assign sub_440_57_n_31 = ~({in1[10]} | {in1[11]});
 assign sub_440_57_n_30 = ~({in1[18]} | {in1[19]});
 assign sub_440_57_n_29 = ~({in1[14]} | {in1[15]});
 assign sub_440_57_n_28 = ~({in1[12]} | {in1[13]});
 assign sub_440_57_n_37 = ~(sub_440_57_n_15 & R_25_6_);
 assign sub_440_57_n_36 = ~(R_25_5_ & ~{in1[6]});
 assign sub_440_57_n_35 = ~(R_25_4_ | ~{in1[5]});
 assign sub_440_57_n_11 = ~(R_25_4_ & ~{in1[5]});
 assign sub_440_57_n_34 = ~(sub_440_57_n_14 & R_25_1_);
 assign sub_440_57_n_32 = ~(R_25_2_ | ~{in1[3]});
 assign sub_440_57_n_25 = ~sub_440_57_n_2;
 assign sub_440_57_n_20 = ~({in1[20]} | {in1[21]});
 assign sub_440_57_n_19 = ~({in1[8]} | {in1[9]});
 assign sub_440_57_n_18 = ~({in1[16]} | {in1[17]});
 assign sub_440_57_n_17 = ~({in1[22]} | {in1[23]});
 assign sub_440_57_n_27 = ~(sub_440_57_n_16 & ~sub_440_57_n_14);
 assign sub_440_57_n_26 = ~(R_25_0_ & ~{in1[1]});
 assign sub_440_57_n_24 = ~(R_25_3_ | ~{in1[4]});
 assign sub_440_57_n_23 = ~(R_25_6_ | ~{in1[7]});
 assign sub_440_57_n_22 = ~(R_25_5_ | ~{in1[6]});
 assign sub_440_57_n_21 = ~({in2[24]} | ~{in1[0]});
 assign sub_440_57_n_16 = ~R_25_1_;
 assign sub_440_57_n_15 = ~{in1[7]};
 assign sub_440_57_n_14 = ~{in1[2]};
 assign sub_440_57_n_10 = ~({in1[4]} & ~R_25_3_);
 assign sub_440_57_n_9 = ~(sub_440_57_n_23 | ~sub_440_57_n_37);
 assign sub_440_57_n_8 = ~(sub_440_57_n_22 | ~sub_440_57_n_36);
 assign sub_440_57_n_7 = ~(sub_440_57_n_21 | ~sub_440_57_n_4);
 assign sub_440_57_n_6 = ~(sub_440_57_n_2 & ~sub_440_57_n_24);
 assign sub_440_57_n_5 = (R_25_6_ | sub_440_57_n_15);
 assign sub_440_57_n_4 = ~({in1[1]} & ~R_25_0_);
 assign sub_440_57_n_3 = ~({in1[6]} & ~R_25_5_);
 assign sub_440_57_n_2 = ~(R_25_3_ & ~{in1[4]});
 assign sub_440_57_n_1 = ~({in1[5]} & ~R_25_4_);
 assign sub_440_57_n_0 = ~(R_25_2_ & ~{in1[3]});
 assign T_23_7_ = ((sub_470_56_n_66 & sub_470_56_n_3) | ~(sub_470_56_n_66 | sub_470_56_n_3));
 assign T_23_32_ = ~(sub_470_56_n_61 & ~sub_470_56_n_42);
 assign sub_470_56_n_66 = ~(sub_470_56_n_62 & ~sub_470_56_n_24);
 assign T_23_8_ = ~((sub_470_56_n_60 | sub_470_56_n_34) & ~(sub_470_56_n_60 & sub_470_56_n_34));
 assign T_23_6_ = ((sub_470_56_n_59 & sub_470_56_n_8) | ~(sub_470_56_n_59 | sub_470_56_n_8));
 assign T_23_5_ = ~((sub_470_56_n_7 | sub_470_56_n_6) & ~(sub_470_56_n_7 & sub_470_56_n_6));
 assign sub_470_56_n_62 = ~(sub_470_56_n_59 & ~sub_470_56_n_22);
 assign sub_470_56_n_61 = ~(sub_470_56_n_56 & sub_470_56_n_49);
 assign sub_470_56_n_60 = ~(sub_470_56_n_48 & (sub_470_56_n_53 | sub_470_56_n_41));
 assign sub_470_56_n_59 = ~(sub_470_56_n_39 & (~sub_470_56_n_35 | sub_470_56_n_53));
 assign T_23_3_ = ~((sub_470_56_n_54 | sub_470_56_n_9) & ~(sub_470_56_n_54 & sub_470_56_n_9));
 assign T_23_4_ = ((sub_470_56_n_53 & sub_470_56_n_4) | ~(sub_470_56_n_53 | sub_470_56_n_4));
 assign sub_470_56_n_56 = ~(sub_470_56_n_55 | ~sub_470_56_n_10);
 assign sub_470_56_n_55 = ~(sub_470_56_n_44 | (sub_470_56_n_41 | sub_470_56_n_53));
 assign sub_470_56_n_54 = ~(sub_470_56_n_0 & (sub_470_56_n_46 | sub_470_56_n_19));
 assign sub_470_56_n_53 = ~(sub_470_56_n_51 | sub_470_56_n_37);
 assign T_23_2_ = ~((sub_470_56_n_50 | sub_470_56_n_5) & ~(sub_470_56_n_50 & sub_470_56_n_5));
 assign sub_470_56_n_51 = ~(sub_470_56_n_19 | (sub_470_56_n_23 | sub_470_56_n_46));
 assign sub_470_56_n_50 = ~sub_470_56_n_46;
 assign sub_470_56_n_49 = ~(sub_470_56_n_47 & ~sub_470_56_n_44);
 assign sub_470_56_n_48 = ~sub_470_56_n_47;
 assign sub_470_56_n_47 = ~(sub_470_56_n_43 & ~sub_470_56_n_36);
 assign sub_470_56_n_46 = ~((n_1019 & R_24_0_) | ((R_24_0_ & sub_470_56_n_15) | (sub_470_56_n_15 & n_1019)));
 assign T_23_1_ = ~(R_24_0_ ^ (n_1349 ^ n_1019));
 assign sub_470_56_n_44 = ~(sub_470_56_n_40 & sub_470_56_n_1);
 assign sub_470_56_n_43 = ~(sub_470_56_n_38 & sub_470_56_n_33);
 assign sub_470_56_n_42 = ~(sub_470_56_n_31 & (sub_470_56_n_32 & (sub_470_56_n_27 & sub_470_56_n_29)));
 assign sub_470_56_n_41 = ~(sub_470_56_n_35 & sub_470_56_n_33);
 assign sub_470_56_n_40 = ~(n_1344 | (n_1064 | (n_1090 | ~sub_470_56_n_28)));
 assign sub_470_56_n_39 = ~sub_470_56_n_38;
 assign sub_470_56_n_38 = ~(sub_470_56_n_26 & (sub_470_56_n_2 | sub_470_56_n_20));
 assign sub_470_56_n_37 = ~(sub_470_56_n_25 & (sub_470_56_n_0 | sub_470_56_n_23));
 assign sub_470_56_n_36 = ~(sub_470_56_n_21 & (sub_470_56_n_12 | sub_470_56_n_18));
 assign sub_470_56_n_35 = ~(sub_470_56_n_11 | sub_470_56_n_20);
 assign sub_470_56_n_34 = ~(sub_470_56_n_13 & sub_470_56_n_1);
 assign sub_470_56_n_32 = ~(n_1211 | (n_1365 | (n_1176 | n_1291)));
 assign sub_470_56_n_31 = ~(n_1135 | (n_1171 | (n_1030 | n_1301)));
 assign T_23_0_ = ~(sub_470_56_n_17 & (~{in2[23]} | {in1[0]}));
 assign sub_470_56_n_29 = ~(n_1296 | (n_1360 | (n_829 | n_1272)));
 assign sub_470_56_n_28 = ~(n_1161 | (n_1025 | (n_1258 | n_1181)));
 assign sub_470_56_n_27 = ~(n_1058 | (n_1370 | (n_1085 | n_1241)));
 assign sub_470_56_n_33 = ~(sub_470_56_n_22 | sub_470_56_n_18);
 assign sub_470_56_n_24 = ~sub_470_56_n_12;
 assign sub_470_56_n_13 = ~(sub_470_56_n_16 & R_24_7_);
 assign sub_470_56_n_26 = ~(R_24_4_ & ~n_1048);
 assign sub_470_56_n_25 = ~(R_24_2_ & ~n_1112);
 assign sub_470_56_n_12 = ~(R_24_5_ & ~n_1095);
 assign sub_470_56_n_23 = ~(R_24_2_ | ~n_1112);
 assign sub_470_56_n_22 = ~(R_24_5_ | ~n_1095);
 assign sub_470_56_n_21 = ~(R_24_6_ & ~n_1166);
 assign sub_470_56_n_11 = ~(R_24_3_ | ~n_1339);
 assign sub_470_56_n_20 = ~(R_24_4_ | ~n_1048);
 assign sub_470_56_n_19 = ~(R_24_1_ | ~n_1100);
 assign sub_470_56_n_18 = ~(R_24_6_ | ~n_1166);
 assign sub_470_56_n_17 = ~({in1[0]} & ~{in2[23]});
 assign sub_470_56_n_16 = ~n_1216;
 assign sub_470_56_n_15 = ~n_1349;
 assign sub_470_56_n_10 = ~(sub_470_56_n_40 & ~sub_470_56_n_13);
 assign sub_470_56_n_9 = ~(sub_470_56_n_25 & ~sub_470_56_n_23);
 assign sub_470_56_n_8 = ~(sub_470_56_n_12 & ~sub_470_56_n_22);
 assign sub_470_56_n_7 = ~(sub_470_56_n_2 & (sub_470_56_n_11 | sub_470_56_n_53));
 assign sub_470_56_n_6 = ~(sub_470_56_n_26 & ~sub_470_56_n_20);
 assign sub_470_56_n_5 = ~(sub_470_56_n_0 & ~sub_470_56_n_19);
 assign sub_470_56_n_4 = ~(sub_470_56_n_11 | ~sub_470_56_n_2);
 assign sub_470_56_n_3 = ~(sub_470_56_n_21 & ~sub_470_56_n_18);
 assign sub_470_56_n_2 = ~(R_24_3_ & ~n_1339);
 assign sub_470_56_n_1 = (R_24_7_ | sub_470_56_n_16);
 assign sub_470_56_n_0 = ~(R_24_1_ & ~n_1100);
 assign T_22_9_ = ((sub_500_55_n_85 & sub_500_55_n_13) | ~(sub_500_55_n_85 | sub_500_55_n_13));
 assign T_22_7_ = ((sub_500_55_n_8 & ~sub_500_55_n_81) | (sub_500_55_n_39 & sub_500_55_n_81));
 assign sub_500_55_n_85 = ~(sub_500_55_n_28 & (~sub_500_55_n_6 | sub_500_55_n_79));
 assign T_22_5_ = ((sub_500_55_n_7 & ~sub_500_55_n_77) | (sub_500_55_n_52 & sub_500_55_n_77));
 assign T_22_8_ = ((sub_500_55_n_80 & sub_500_55_n_48) | ~(sub_500_55_n_80 | sub_500_55_n_48));
 assign T_22_32_ = ~(sub_500_55_n_78 & ~sub_500_55_n_18);
 assign sub_500_55_n_81 = ~(sub_500_55_n_3 | (~sub_500_55_n_37 & sub_500_55_n_75));
 assign sub_500_55_n_80 = ~sub_500_55_n_79;
 assign sub_500_55_n_79 = ~(sub_500_55_n_14 | (~sub_500_55_n_60 & sub_500_55_n_73));
 assign sub_500_55_n_78 = ~(sub_500_55_n_70 & sub_500_55_n_74);
 assign sub_500_55_n_77 = ~(sub_500_55_n_0 | (~sub_500_55_n_29 & sub_500_55_n_73));
 assign T_22_4_ = ~((sub_500_55_n_73 | sub_500_55_n_11) & ~(sub_500_55_n_73 & sub_500_55_n_11));
 assign sub_500_55_n_75 = ~(sub_500_55_n_57 & (sub_500_55_n_68 | sub_500_55_n_55));
 assign sub_500_55_n_74 = ~(sub_500_55_n_73 & ~sub_500_55_n_60);
 assign sub_500_55_n_73 = ~(sub_500_55_n_69 & ~sub_500_55_n_56);
 assign sub_500_55_n_72 = ~(sub_500_55_n_32 | (~sub_500_55_n_34 & sub_500_55_n_66));
 assign T_22_2_ = ~((sub_500_55_n_66 | sub_500_55_n_10) & ~(sub_500_55_n_66 & sub_500_55_n_10));
 assign sub_500_55_n_70 = ~(sub_500_55_n_14 | ~sub_500_55_n_67);
 assign sub_500_55_n_69 = ~(sub_500_55_n_64 & (sub_500_55_n_25 & sub_500_55_n_51));
 assign sub_500_55_n_68 = ~(sub_500_55_n_49 | (sub_500_55_n_64 & sub_500_55_n_51));
 assign sub_500_55_n_67 = ~(sub_500_55_n_63 & sub_500_55_n_41);
 assign sub_500_55_n_66 = ~(sub_500_55_n_2 & (sub_500_55_n_23 | sub_500_55_n_33));
 assign T_22_1_ = ~((sub_500_55_n_9 | sub_500_55_n_61) & ~(sub_500_55_n_9 & sub_500_55_n_61));
 assign sub_500_55_n_64 = ~(sub_500_55_n_23 & sub_500_55_n_2);
 assign sub_500_55_n_63 = ~(sub_500_55_n_59 | sub_500_55_n_38);
 assign sub_500_55_n_62 = (sub_500_55_n_45 & (sub_500_55_n_42 & (sub_500_55_n_44 & sub_500_55_n_40)));
 assign sub_500_55_n_61 = ~sub_500_55_n_23;
 assign sub_500_55_n_60 = ~(sub_500_55_n_53 & sub_500_55_n_47);
 assign sub_500_55_n_59 = (n_1181 | (n_1090 | sub_500_55_n_43));
 assign sub_500_55_n_58 = ~(sub_500_55_n_30 | (sub_500_55_n_3 & sub_500_55_n_1));
 assign sub_500_55_n_57 = ~(sub_500_55_n_5 | (sub_500_55_n_0 & sub_500_55_n_36));
 assign sub_500_55_n_56 = ~(sub_500_55_n_24 & (sub_500_55_n_4 | sub_500_55_n_26));
 assign sub_500_55_n_55 = ~(sub_500_55_n_50 & sub_500_55_n_53);
 assign sub_500_55_n_52 = ~sub_500_55_n_7;
 assign sub_500_55_n_50 = ~(sub_500_55_n_26 & sub_500_55_n_24);
 assign sub_500_55_n_49 = ~(sub_500_55_n_4 & sub_500_55_n_24);
 assign sub_500_55_n_54 = ~(sub_500_55_n_24 & sub_500_55_n_25);
 assign sub_500_55_n_53 = ~(sub_500_55_n_29 | sub_500_55_n_35);
 assign sub_500_55_n_51 = ~(sub_500_55_n_33 | sub_500_55_n_34);
 assign T_22_0_ = (sub_500_55_n_23 | (n_1323 & n_1057));
 assign sub_500_55_n_45 = ~(n_1135 | (n_1171 | (n_1030 | n_1301)));
 assign sub_500_55_n_44 = ~(n_1058 | (n_1370 | (n_1085 | n_1241)));
 assign sub_500_55_n_43 = (n_1344 | (n_1064 | (n_1025 | n_1258)));
 assign sub_500_55_n_42 = ~(n_1211 | (n_1365 | (n_1176 | n_1291)));
 assign sub_500_55_n_41 = ~(sub_500_55_n_28 & sub_500_55_n_31);
 assign sub_500_55_n_40 = ~(n_1296 | (n_1360 | (n_829 | n_1272)));
 assign sub_500_55_n_48 = ~(sub_500_55_n_28 & sub_500_55_n_6);
 assign sub_500_55_n_47 = ~(sub_500_55_n_37 | sub_500_55_n_27);
 assign sub_500_55_n_39 = ~(sub_500_55_n_30 | sub_500_55_n_27);
 assign sub_500_55_n_36 = ~sub_500_55_n_35;
 assign sub_500_55_n_32 = ~sub_500_55_n_4;
 assign sub_500_55_n_38 = ~(R_23_8_ | ~n_1161);
 assign sub_500_55_n_37 = ~(R_23_5_ | ~n_1095);
 assign sub_500_55_n_35 = ~(R_23_4_ | ~n_1048);
 assign sub_500_55_n_34 = ~(R_23_1_ | ~n_1100);
 assign sub_500_55_n_33 = ~(R_23_0_ | ~n_1349);
 assign sub_500_55_n_25 = ~sub_500_55_n_26;
 assign sub_500_55_n_31 = ~(R_23_8_ & ~n_1161);
 assign sub_500_55_n_30 = ~(n_1166 | sub_500_55_n_21);
 assign sub_500_55_n_29 = ~(R_23_3_ | ~n_1339);
 assign sub_500_55_n_28 = ~(sub_500_55_n_22 & R_23_7_);
 assign sub_500_55_n_27 = ~(R_23_6_ | ~n_1166);
 assign sub_500_55_n_26 = ~(R_23_2_ | ~n_1112);
 assign sub_500_55_n_24 = ~(R_23_2_ & ~n_1112);
 assign sub_500_55_n_23 = ~(n_1057 | n_1323);
 assign sub_500_55_n_22 = ~n_1216;
 assign sub_500_55_n_21 = ~R_23_6_;
 assign sub_500_55_n_20 = ~{in1[0]};
 assign sub_500_55_n_18 = ~(sub_500_55_n_62 & (~sub_500_55_n_67 | sub_500_55_n_17));
 assign sub_500_55_n_17 = (sub_500_55_n_63 & sub_500_55_n_6);
 assign T_22_3_ = (sub_500_55_n_72 ^ sub_500_55_n_54);
 assign T_22_6_ = ~(sub_500_55_n_75 ^ sub_500_55_n_12);
 assign sub_500_55_n_14 = ~(sub_500_55_n_58 & (~sub_500_55_n_47 | sub_500_55_n_57));
 assign sub_500_55_n_13 = ~(sub_500_55_n_31 & ~sub_500_55_n_38);
 assign sub_500_55_n_12 = (sub_500_55_n_3 | sub_500_55_n_37);
 assign sub_500_55_n_11 = (sub_500_55_n_0 | sub_500_55_n_29);
 assign sub_500_55_n_10 = ~(sub_500_55_n_4 & ~sub_500_55_n_34);
 assign sub_500_55_n_9 = ~(sub_500_55_n_2 & ~sub_500_55_n_33);
 assign sub_500_55_n_8 = ~(sub_500_55_n_1 & ~sub_500_55_n_30);
 assign sub_500_55_n_7 = ~(sub_500_55_n_36 & ~sub_500_55_n_5);
 assign sub_500_55_n_6 = (R_23_7_ | sub_500_55_n_22);
 assign sub_500_55_n_5 = ~(n_1048 | ~R_23_4_);
 assign sub_500_55_n_4 = ~(R_23_1_ & ~n_1100);
 assign sub_500_55_n_3 = ~(n_1095 | ~R_23_5_);
 assign sub_500_55_n_2 = ~(R_23_0_ & ~n_1349);
 assign sub_500_55_n_1 = ~(sub_500_55_n_21 & n_1166);
 assign sub_500_55_n_0 = ~(n_1339 | ~R_23_3_);
 assign T_21_10_ = ((sub_530_54_n_88 & sub_530_54_n_8) | ~(sub_530_54_n_88 | sub_530_54_n_8));
 assign T_21_7_ = ~((sub_530_54_n_89 | sub_530_54_n_56) & ~(sub_530_54_n_89 & sub_530_54_n_56));
 assign T_21_9_ = ((sub_530_54_n_87 & sub_530_54_n_6) | ~(sub_530_54_n_87 | sub_530_54_n_6));
 assign sub_530_54_n_89 = ~(sub_530_54_n_2 | (~sub_530_54_n_38 & sub_530_54_n_81));
 assign sub_530_54_n_88 = ~(sub_530_54_n_59 & (~sub_530_54_n_45 | sub_530_54_n_16));
 assign sub_530_54_n_87 = ~(sub_530_54_n_0 & (~sub_530_54_n_32 | sub_530_54_n_16));
 assign T_21_8_ = ((sub_530_54_n_21 & sub_530_54_n_52) | ~(sub_530_54_n_21 | sub_530_54_n_52));
 assign T_21_6_ = ((sub_530_54_n_81 & sub_530_54_n_13) | ~(sub_530_54_n_81 | sub_530_54_n_13));
 assign T_21_5_ = ((sub_530_54_n_11 & sub_530_54_n_12) | ~(sub_530_54_n_11 | sub_530_54_n_12));
 assign T_21_32_ = ~(sub_530_54_n_82 & ~sub_530_54_n_71);
 assign sub_530_54_n_21 = ~sub_530_54_n_16;
 assign sub_530_54_n_82 = ~(sub_530_54_n_70 & sub_530_54_n_79);
 assign sub_530_54_n_81 = ~(sub_530_54_n_57 & (~sub_530_54_n_53 | sub_530_54_n_77));
 assign T_21_4_ = ~((sub_530_54_n_77 | sub_530_54_n_7) & ~(sub_530_54_n_77 & sub_530_54_n_7));
 assign sub_530_54_n_79 = ~(sub_530_54_n_76 & ~sub_530_54_n_62);
 assign sub_530_54_n_78 = ~(sub_530_54_n_18 & (sub_530_54_n_72 | sub_530_54_n_36));
 assign sub_530_54_n_77 = ~sub_530_54_n_76;
 assign sub_530_54_n_76 = ~(sub_530_54_n_74 & sub_530_54_n_61);
 assign T_21_2_ = ~((sub_530_54_n_73 | sub_530_54_n_10) & ~(sub_530_54_n_73 & sub_530_54_n_10));
 assign sub_530_54_n_74 = ~(sub_530_54_n_67 & sub_530_54_n_50);
 assign sub_530_54_n_73 = ~sub_530_54_n_72;
 assign sub_530_54_n_72 = ~sub_530_54_n_67;
 assign sub_530_54_n_71 = ~(sub_530_54_n_69 & (sub_530_54_n_55 | (sub_530_54_n_60 & sub_530_54_n_51)));
 assign sub_530_54_n_70 = ~(sub_530_54_n_68 | ~sub_530_54_n_65);
 assign sub_530_54_n_69 = (sub_530_54_n_44 & (sub_530_54_n_42 & (sub_530_54_n_41 & sub_530_54_n_63)));
 assign sub_530_54_n_68 = ~(sub_530_54_n_14 & (~sub_530_54_n_48 | sub_530_54_n_57));
 assign sub_530_54_n_67 = ~(sub_530_54_n_1 & (sub_530_54_n_26 | sub_530_54_n_30));
 assign T_21_1_ = ((sub_530_54_n_9 & sub_530_54_n_64) | ~(sub_530_54_n_9 | sub_530_54_n_64));
 assign sub_530_54_n_65 = ~(sub_530_54_n_58 | sub_530_54_n_55);
 assign sub_530_54_n_64 = ~sub_530_54_n_26;
 assign sub_530_54_n_63 = (sub_530_54_n_46 & sub_530_54_n_43);
 assign sub_530_54_n_62 = ~(sub_530_54_n_53 & sub_530_54_n_48);
 assign sub_530_54_n_61 = ~(sub_530_54_n_40 | (sub_530_54_n_35 & sub_530_54_n_34));
 assign sub_530_54_n_60 = ~(sub_530_54_n_27 | (sub_530_54_n_31 & sub_530_54_n_3));
 assign sub_530_54_n_59 = ~sub_530_54_n_58;
 assign sub_530_54_n_58 = ~(sub_530_54_n_3 & (sub_530_54_n_0 | sub_530_54_n_25));
 assign sub_530_54_n_57 = ~(sub_530_54_n_49 | ~sub_530_54_n_4);
 assign sub_530_54_n_51 = ~(sub_530_54_n_28 | ~sub_530_54_n_23);
 assign sub_530_54_n_50 = ~(sub_530_54_n_36 | sub_530_54_n_33);
 assign sub_530_54_n_49 = ~(sub_530_54_n_5 | sub_530_54_n_37);
 assign sub_530_54_n_56 = ~(sub_530_54_n_17 | sub_530_54_n_39);
 assign sub_530_54_n_55 = ~(sub_530_54_n_29 | ~sub_530_54_n_23);
 assign sub_530_54_n_54 = ~(sub_530_54_n_20 & sub_530_54_n_34);
 assign sub_530_54_n_53 = ~(sub_530_54_n_19 | sub_530_54_n_37);
 assign sub_530_54_n_52 = ~(sub_530_54_n_0 & sub_530_54_n_32);
 assign T_21_0_ = (sub_530_54_n_26 | (n_1322 & n_1018));
 assign sub_530_54_n_46 = ~(n_1211 | (n_1365 | (n_1176 | n_1291)));
 assign sub_530_54_n_45 = ~(sub_530_54_n_31 | sub_530_54_n_27);
 assign sub_530_54_n_44 = ~(n_1025 | (n_1258 | (n_1181 | n_1090)));
 assign sub_530_54_n_43 = ~(n_1058 | (n_1370 | (n_1085 | n_1241)));
 assign sub_530_54_n_42 = ~(n_1135 | (n_1171 | (n_1030 | n_1301)));
 assign sub_530_54_n_41 = ~(n_1296 | (n_1360 | (n_829 | n_1272)));
 assign sub_530_54_n_48 = ~(sub_530_54_n_38 | sub_530_54_n_39);
 assign sub_530_54_n_40 = ~sub_530_54_n_20;
 assign sub_530_54_n_35 = ~sub_530_54_n_18;
 assign sub_530_54_n_34 = ~sub_530_54_n_33;
 assign sub_530_54_n_32 = ~sub_530_54_n_31;
 assign sub_530_54_n_20 = ~(R_22_2_ & ~n_1112);
 assign sub_530_54_n_39 = ~(R_22_6_ | ~n_1166);
 assign sub_530_54_n_38 = ~(R_22_5_ | ~n_1095);
 assign sub_530_54_n_37 = ~(R_22_4_ | ~n_1048);
 assign sub_530_54_n_19 = ~(R_22_3_ | ~n_1339);
 assign sub_530_54_n_36 = ~(R_22_1_ | ~n_1100);
 assign sub_530_54_n_18 = ~(R_22_1_ & ~n_1100);
 assign sub_530_54_n_33 = ~(R_22_2_ | ~n_1112);
 assign sub_530_54_n_31 = ~(R_22_7_ | ~n_1216);
 assign sub_530_54_n_30 = ~(R_22_0_ | ~n_1349);
 assign sub_530_54_n_29 = ~(R_22_9_ & ~n_1344);
 assign sub_530_54_n_28 = ~(R_22_9_ | ~n_1344);
 assign sub_530_54_n_25 = ~(R_22_8_ | ~n_1161);
 assign sub_530_54_n_27 = ~(R_22_8_ | ~n_1161);
 assign sub_530_54_n_26 = ~(n_1018 | n_1322);
 assign sub_530_54_n_24 = ~{in1[0]};
 assign sub_530_54_n_23 = ~n_1064;
 assign sub_530_54_n_17 = ~(n_1166 | ~R_22_6_);
 assign sub_530_54_n_16 = ~(sub_530_54_n_68 | ~sub_530_54_n_79);
 assign T_21_3_ = ~(sub_530_54_n_78 ^ sub_530_54_n_54);
 assign sub_530_54_n_14 = ~(sub_530_54_n_17 | (~sub_530_54_n_39 & sub_530_54_n_2));
 assign sub_530_54_n_13 = (sub_530_54_n_2 | sub_530_54_n_38);
 assign sub_530_54_n_12 = ~(sub_530_54_n_4 & ~sub_530_54_n_37);
 assign sub_530_54_n_11 = ~(sub_530_54_n_5 & (sub_530_54_n_19 | sub_530_54_n_77));
 assign sub_530_54_n_10 = ~(sub_530_54_n_18 & ~sub_530_54_n_36);
 assign sub_530_54_n_9 = ~(sub_530_54_n_1 & ~sub_530_54_n_30);
 assign sub_530_54_n_8 = ~(sub_530_54_n_29 & ~sub_530_54_n_28);
 assign sub_530_54_n_7 = ~(sub_530_54_n_19 | ~sub_530_54_n_5);
 assign sub_530_54_n_6 = ~(sub_530_54_n_3 & ~sub_530_54_n_27);
 assign sub_530_54_n_5 = ~(R_22_3_ & ~n_1339);
 assign sub_530_54_n_4 = ~(R_22_4_ & ~n_1048);
 assign sub_530_54_n_3 = ~(R_22_8_ & ~n_1161);
 assign sub_530_54_n_2 = ~(n_1095 | ~R_22_5_);
 assign sub_530_54_n_1 = ~(R_22_0_ & ~n_1349);
 assign sub_530_54_n_0 = ~(R_22_7_ & ~n_1216);
 assign T_20_11_ = ((sub_560_53_n_103 & sub_560_53_n_14) | ~(sub_560_53_n_103 | sub_560_53_n_14));
 assign sub_560_53_n_103 = ~(sub_560_53_n_9 & (~sub_560_53_n_41 | sub_560_53_n_95));
 assign T_20_10_ = ~((sub_560_53_n_95 | sub_560_53_n_11) & ~(sub_560_53_n_95 & sub_560_53_n_11));
 assign T_20_9_ = ~((sub_560_53_n_97 | sub_560_53_n_13) & ~(sub_560_53_n_97 & sub_560_53_n_13));
 assign T_20_7_ = ~((sub_560_53_n_96 | sub_560_53_n_15) & ~(sub_560_53_n_96 & sub_560_53_n_15));
 assign T_20_32_ = ~(sub_560_53_n_98 & ~sub_560_53_n_68);
 assign sub_560_53_n_98 = ~(sub_560_53_n_91 & ~sub_560_53_n_79);
 assign sub_560_53_n_97 = ~(sub_560_53_n_39 & (~sub_560_53_n_10 | sub_560_53_n_89));
 assign sub_560_53_n_96 = ~(sub_560_53_n_5 | (sub_560_53_n_84 & sub_560_53_n_4));
 assign sub_560_53_n_95 = ~(sub_560_53_n_60 | (~sub_560_53_n_48 & sub_560_53_n_88));
 assign T_20_8_ = ((sub_560_53_n_89 & sub_560_53_n_19) | ~(sub_560_53_n_89 | sub_560_53_n_19));
 assign T_20_6_ = ((sub_560_53_n_85 & sub_560_53_n_17) | ~(sub_560_53_n_85 | sub_560_53_n_17));
 assign T_20_5_ = ((sub_560_53_n_87 & sub_560_53_n_12) | ~(sub_560_53_n_87 | sub_560_53_n_12));
 assign sub_560_53_n_91 = ~(sub_560_53_n_88 & ~sub_560_53_n_70);
 assign T_20_3_ = ((sub_560_53_n_82 & sub_560_53_n_50) | ~(sub_560_53_n_82 | sub_560_53_n_50));
 assign sub_560_53_n_89 = ~sub_560_53_n_88;
 assign sub_560_53_n_88 = ~(sub_560_53_n_81 & ~(sub_560_53_n_78 & sub_560_53_n_55));
 assign sub_560_53_n_87 = ~(sub_560_53_n_2 | (sub_560_53_n_20 & sub_560_53_n_8));
 assign T_20_4_ = ~((sub_560_53_n_20 | sub_560_53_n_16) & ~(sub_560_53_n_20 & sub_560_53_n_16));
 assign sub_560_53_n_85 = ~sub_560_53_n_84;
 assign sub_560_53_n_84 = ~(sub_560_53_n_83 & ~sub_560_53_n_64);
 assign sub_560_53_n_83 = ~(sub_560_53_n_20 & ~sub_560_53_n_56);
 assign sub_560_53_n_82 = ~(sub_560_53_n_35 & (~sub_560_53_n_38 | sub_560_53_n_76));
 assign sub_560_53_n_81 = ~(sub_560_53_n_69 | (sub_560_53_n_75 & sub_560_53_n_63));
 assign T_20_2_ = ((sub_560_53_n_77 & sub_560_53_n_58) | ~(sub_560_53_n_77 | sub_560_53_n_58));
 assign sub_560_53_n_79 = ~(sub_560_53_n_51 | (sub_560_53_n_73 & sub_560_53_n_62));
 assign sub_560_53_n_78 = ~(sub_560_53_n_37 & (sub_560_53_n_71 | sub_560_53_n_56));
 assign sub_560_53_n_77 = ~sub_560_53_n_76;
 assign sub_560_53_n_76 = ~(sub_560_53_n_18 | ~sub_560_53_n_31);
 assign sub_560_53_n_75 = ~(sub_560_53_n_59 | ~sub_560_53_n_72);
 assign T_20_1_ = ((sub_560_53_n_57 & sub_560_53_n_66) | ~(sub_560_53_n_57 | sub_560_53_n_66));
 assign sub_560_53_n_73 = ~(sub_560_53_n_60 & sub_560_53_n_49);
 assign sub_560_53_n_72 = ~(sub_560_53_n_30 & sub_560_53_n_31);
 assign sub_560_53_n_71 = ~(sub_560_53_n_67 | (sub_560_53_n_29 & sub_560_53_n_0));
 assign sub_560_53_n_70 = ~(sub_560_53_n_65 & sub_560_53_n_49);
 assign sub_560_53_n_69 = ~(sub_560_53_n_61 & (sub_560_53_n_52 | sub_560_53_n_54));
 assign sub_560_53_n_68 = ~(sub_560_53_n_46 & (sub_560_53_n_44 & (sub_560_53_n_45 & sub_560_53_n_43)));
 assign sub_560_53_n_67 = ~sub_560_53_n_42;
 assign sub_560_53_n_66 = ~sub_560_53_n_30;
 assign sub_560_53_n_65 = ~(sub_560_53_n_51 | sub_560_53_n_48);
 assign sub_560_53_n_64 = ~(sub_560_53_n_52 & ~sub_560_53_n_21);
 assign sub_560_53_n_63 = ~(sub_560_53_n_56 | sub_560_53_n_54);
 assign sub_560_53_n_62 = ~(sub_560_53_n_53 | ~sub_560_53_n_7);
 assign sub_560_53_n_61 = ~(sub_560_53_n_36 | (sub_560_53_n_5 & sub_560_53_n_3));
 assign sub_560_53_n_60 = ~(sub_560_53_n_34 & (sub_560_53_n_39 | sub_560_53_n_32));
 assign sub_560_53_n_59 = ~(sub_560_53_n_38 & (sub_560_53_n_0 & sub_560_53_n_6));
 assign sub_560_53_n_55 = ~sub_560_53_n_54;
 assign sub_560_53_n_53 = ~(sub_560_53_n_9 | sub_560_53_n_33);
 assign sub_560_53_n_58 = ~(sub_560_53_n_35 & sub_560_53_n_38);
 assign sub_560_53_n_57 = ~(sub_560_53_n_31 & sub_560_53_n_6);
 assign sub_560_53_n_56 = ~(sub_560_53_n_8 & sub_560_53_n_1);
 assign sub_560_53_n_54 = ~(sub_560_53_n_4 & sub_560_53_n_3);
 assign T_20_0_ = (sub_560_53_n_30 | (n_1321 & n_1109));
 assign sub_560_53_n_46 = ~(n_1135 | (n_1171 | (n_1030 | n_1301)));
 assign sub_560_53_n_45 = ~(n_1058 | (n_1370 | (n_1085 | n_1241)));
 assign sub_560_53_n_44 = ~(n_1211 | (n_1365 | (n_1176 | n_1291)));
 assign sub_560_53_n_43 = ~(n_1296 | (n_1360 | (n_829 | n_1272)));
 assign sub_560_53_n_52 = ~(sub_560_53_n_2 & sub_560_53_n_1);
 assign sub_560_53_n_51 = (n_1025 | (n_1258 | (n_1181 | n_1090)));
 assign sub_560_53_n_50 = ~(sub_560_53_n_42 & (~n_1112 | R_21_2_));
 assign sub_560_53_n_49 = ~(sub_560_53_n_40 | sub_560_53_n_33);
 assign sub_560_53_n_48 = ~(sub_560_53_n_10 & ~sub_560_53_n_32);
 assign sub_560_53_n_41 = ~sub_560_53_n_40;
 assign sub_560_53_n_37 = ~sub_560_53_n_21;
 assign sub_560_53_n_42 = ~(R_21_2_ & ~n_1112);
 assign sub_560_53_n_40 = ~(R_21_9_ | ~n_1344);
 assign sub_560_53_n_39 = ~(R_21_7_ & ~n_1216);
 assign sub_560_53_n_38 = ~(sub_560_53_n_28 & ~sub_560_53_n_23);
 assign sub_560_53_n_21 = ~(n_1048 | sub_560_53_n_27);
 assign sub_560_53_n_29 = ~(n_1100 | sub_560_53_n_28);
 assign sub_560_53_n_36 = ~(n_1166 | sub_560_53_n_24);
 assign sub_560_53_n_35 = ~(sub_560_53_n_23 & R_21_1_);
 assign sub_560_53_n_34 = ~(R_21_8_ & ~n_1161);
 assign sub_560_53_n_33 = ~(R_21_10_ | ~n_1064);
 assign sub_560_53_n_32 = ~(R_21_8_ | ~n_1161);
 assign sub_560_53_n_31 = ~(sub_560_53_n_26 & R_21_0_);
 assign sub_560_53_n_30 = ~(n_1109 | n_1321);
 assign sub_560_53_n_28 = ~R_21_1_;
 assign sub_560_53_n_27 = ~R_21_4_;
 assign sub_560_53_n_26 = ~n_1349;
 assign sub_560_53_n_25 = ~{in1[0]};
 assign sub_560_53_n_24 = ~R_21_6_;
 assign sub_560_53_n_23 = ~n_1100;
 assign sub_560_53_n_20 = ~(sub_560_53_n_71 & ~sub_560_53_n_75);
 assign sub_560_53_n_19 = (sub_560_53_n_39 & sub_560_53_n_10);
 assign sub_560_53_n_18 = ~(sub_560_53_n_30 | ~sub_560_53_n_6);
 assign sub_560_53_n_17 = ~(sub_560_53_n_5 | ~sub_560_53_n_4);
 assign sub_560_53_n_16 = ~(sub_560_53_n_8 & ~sub_560_53_n_2);
 assign sub_560_53_n_15 = ~(sub_560_53_n_36 | ~sub_560_53_n_3);
 assign sub_560_53_n_14 = ~(sub_560_53_n_7 & ~sub_560_53_n_33);
 assign sub_560_53_n_13 = ~(sub_560_53_n_34 & ~sub_560_53_n_32);
 assign sub_560_53_n_12 = ~(sub_560_53_n_21 | ~sub_560_53_n_1);
 assign sub_560_53_n_11 = ~(sub_560_53_n_40 | ~sub_560_53_n_9);
 assign sub_560_53_n_10 = ~(n_1216 & ~R_21_7_);
 assign sub_560_53_n_9 = ~(R_21_9_ & ~n_1344);
 assign sub_560_53_n_8 = ~(n_1339 & ~R_21_3_);
 assign sub_560_53_n_7 = ~(R_21_10_ & ~n_1064);
 assign sub_560_53_n_6 = (R_21_0_ | sub_560_53_n_26);
 assign sub_560_53_n_5 = ~(n_1095 | ~R_21_5_);
 assign sub_560_53_n_4 = ~(n_1095 & ~R_21_5_);
 assign sub_560_53_n_3 = ~(sub_560_53_n_24 & n_1166);
 assign sub_560_53_n_2 = ~(n_1339 | ~R_21_3_);
 assign sub_560_53_n_1 = ~(sub_560_53_n_27 & n_1048);
 assign sub_560_53_n_0 = ~(n_1112 & ~R_21_2_);
 assign T_19_12_ = ((sub_590_52_n_105 & sub_590_52_n_10) | ~(sub_590_52_n_105 | sub_590_52_n_10));
 assign T_19_9_ = ((sub_590_52_n_104 & sub_590_52_n_15) | ~(sub_590_52_n_104 | sub_590_52_n_15));
 assign T_19_11_ = ~((sub_590_52_n_101 | sub_590_52_n_16) & ~(sub_590_52_n_101 & sub_590_52_n_16));
 assign T_19_7_ = ((sub_590_52_n_100 & sub_590_52_n_66) | ~(sub_590_52_n_100 | sub_590_52_n_66));
 assign sub_590_52_n_105 = ~(sub_590_52_n_81 | (~sub_590_52_n_74 & sub_590_52_n_97));
 assign sub_590_52_n_104 = ~(sub_590_52_n_43 | (~sub_590_52_n_46 & sub_590_52_n_97));
 assign T_19_8_ = ~((sub_590_52_n_97 | sub_590_52_n_14) & ~(sub_590_52_n_97 & sub_590_52_n_14));
 assign T_19_32_ = ~(sub_590_52_n_95 & ~sub_590_52_n_87);
 assign sub_590_52_n_101 = ~(sub_590_52_n_96 | ~sub_590_52_n_8);
 assign sub_590_52_n_100 = ~(sub_590_52_n_35 & (~sub_590_52_n_4 | sub_590_52_n_93));
 assign T_19_10_ = ((sub_590_52_n_22 & sub_590_52_n_11) | ~(sub_590_52_n_22 | sub_590_52_n_11));
 assign T_19_6_ = ((sub_590_52_n_23 & sub_590_52_n_64) | ~(sub_590_52_n_23 | sub_590_52_n_64));
 assign sub_590_52_n_97 = ~(sub_590_52_n_94 & ~sub_590_52_n_82);
 assign sub_590_52_n_96 = ~(sub_590_52_n_22 | ~sub_590_52_n_39);
 assign sub_590_52_n_95 = ~(sub_590_52_n_86 & sub_590_52_n_94);
 assign sub_590_52_n_94 = ~(sub_590_52_n_90 & ~sub_590_52_n_63);
 assign sub_590_52_n_93 = ~(sub_590_52_n_90 | ~sub_590_52_n_70);
 assign sub_590_52_n_92 = ~(sub_590_52_n_1 & (sub_590_52_n_26 | sub_590_52_n_45));
 assign T_19_3_ = ((sub_590_52_n_89 & sub_590_52_n_9) | ~(sub_590_52_n_89 | sub_590_52_n_9));
 assign sub_590_52_n_90 = ~(sub_590_52_n_26 | ~sub_590_52_n_65);
 assign sub_590_52_n_89 = ~(sub_590_52_n_32 | (sub_590_52_n_80 & sub_590_52_n_34));
 assign sub_590_52_n_26 = ~(sub_590_52_n_69 | (sub_590_52_n_80 & sub_590_52_n_54));
 assign T_19_2_ = ~((sub_590_52_n_80 | sub_590_52_n_67) & ~(sub_590_52_n_80 & sub_590_52_n_67));
 assign sub_590_52_n_87 = ~(sub_590_52_n_84 & (sub_590_52_n_81 | sub_590_52_n_21));
 assign sub_590_52_n_86 = ~(sub_590_52_n_82 | (sub_590_52_n_25 | sub_590_52_n_81));
 assign sub_590_52_n_85 = ~(sub_590_52_n_20 & (sub_590_52_n_17 | sub_590_52_n_70));
 assign sub_590_52_n_84 = ~sub_590_52_n_83;
 assign sub_590_52_n_83 = ~(sub_590_52_n_76 & (sub_590_52_n_25 | sub_590_52_n_73));
 assign sub_590_52_n_82 = ~(sub_590_52_n_72 & (sub_590_52_n_70 | sub_590_52_n_63));
 assign sub_590_52_n_81 = ~(sub_590_52_n_78 & ~sub_590_52_n_68);
 assign sub_590_52_n_80 = ~(sub_590_52_n_40 & (sub_590_52_n_31 | sub_590_52_n_30));
 assign T_19_1_ = ~((sub_590_52_n_60 | sub_590_52_n_75) & ~(sub_590_52_n_60 & sub_590_52_n_75));
 assign sub_590_52_n_78 = ~(sub_590_52_n_71 & sub_590_52_n_61);
 assign sub_590_52_n_77 = ~(sub_590_52_n_17 | ~sub_590_52_n_65);
 assign sub_590_52_n_76 = (sub_590_52_n_52 & (sub_590_52_n_57 & (sub_590_52_n_51 & sub_590_52_n_53)));
 assign sub_590_52_n_75 = ~sub_590_52_n_31;
 assign sub_590_52_n_73 = ~(sub_590_52_n_62 | sub_590_52_n_49);
 assign sub_590_52_n_74 = ~(sub_590_52_n_59 & sub_590_52_n_61);
 assign sub_590_52_n_25 = ~(sub_590_52_n_62 | sub_590_52_n_42);
 assign sub_590_52_n_69 = ~(sub_590_52_n_41 & (sub_590_52_n_5 | sub_590_52_n_37));
 assign sub_590_52_n_68 = ~(sub_590_52_n_50 & (sub_590_52_n_8 | sub_590_52_n_38));
 assign sub_590_52_n_72 = ~(sub_590_52_n_56 | ~sub_590_52_n_6);
 assign sub_590_52_n_71 = ~(sub_590_52_n_2 & (sub_590_52_n_7 | sub_590_52_n_36));
 assign sub_590_52_n_70 = ~(sub_590_52_n_55 | ~sub_590_52_n_3);
 assign sub_590_52_n_67 = ~(sub_590_52_n_5 & sub_590_52_n_34);
 assign sub_590_52_n_66 = ~(sub_590_52_n_6 & sub_590_52_n_48);
 assign sub_590_52_n_65 = ~(sub_590_52_n_45 | sub_590_52_n_44);
 assign sub_590_52_n_64 = ~(sub_590_52_n_35 & sub_590_52_n_4);
 assign sub_590_52_n_63 = ~(sub_590_52_n_4 & sub_590_52_n_48);
 assign T_19_0_ = (sub_590_52_n_31 | (n_1320 & n_1024));
 assign sub_590_52_n_57 = ~(n_1211 | (n_1365 | (n_1176 | n_1291)));
 assign sub_590_52_n_56 = ~(sub_590_52_n_35 | sub_590_52_n_47);
 assign sub_590_52_n_55 = ~(sub_590_52_n_1 | sub_590_52_n_44);
 assign sub_590_52_n_54 = ~(sub_590_52_n_33 | sub_590_52_n_37);
 assign sub_590_52_n_53 = ~(n_1296 | (n_1360 | (n_829 | n_1272)));
 assign sub_590_52_n_52 = ~(n_1135 | (n_1171 | (n_1030 | n_1301)));
 assign sub_590_52_n_51 = ~(n_1058 | (n_1370 | (n_1085 | n_1241)));
 assign sub_590_52_n_62 = (n_1181 | (n_1090 | n_1258));
 assign sub_590_52_n_61 = ~(sub_590_52_n_24 | sub_590_52_n_38);
 assign sub_590_52_n_60 = ~(sub_590_52_n_40 & sub_590_52_n_0);
 assign sub_590_52_n_59 = ~(sub_590_52_n_46 | sub_590_52_n_36);
 assign sub_590_52_n_48 = ~sub_590_52_n_47;
 assign sub_590_52_n_43 = ~sub_590_52_n_7;
 assign sub_590_52_n_50 = ~(R_20_10_ & ~n_1064);
 assign sub_590_52_n_49 = ~(R_20_11_ | ~n_1025);
 assign sub_590_52_n_47 = ~(R_20_6_ | ~n_1166);
 assign sub_590_52_n_46 = ~(R_20_7_ | ~n_1216);
 assign sub_590_52_n_45 = ~(R_20_3_ | ~n_1339);
 assign sub_590_52_n_44 = ~(R_20_4_ | ~n_1048);
 assign sub_590_52_n_39 = ~sub_590_52_n_24;
 assign sub_590_52_n_34 = ~sub_590_52_n_33;
 assign sub_590_52_n_32 = ~sub_590_52_n_5;
 assign sub_590_52_n_30 = ~(R_20_0_ | ~n_1349);
 assign sub_590_52_n_42 = ~(R_20_11_ & ~n_1025);
 assign sub_590_52_n_41 = ~(R_20_2_ & ~n_1112);
 assign sub_590_52_n_40 = ~(sub_590_52_n_29 & R_20_0_);
 assign sub_590_52_n_24 = ~(R_20_9_ | ~n_1344);
 assign sub_590_52_n_38 = ~(R_20_10_ | ~n_1064);
 assign sub_590_52_n_37 = ~(R_20_2_ | ~n_1112);
 assign sub_590_52_n_36 = ~(R_20_8_ | ~n_1161);
 assign sub_590_52_n_35 = ~(R_20_5_ & ~n_1095);
 assign sub_590_52_n_33 = ~(R_20_1_ | ~n_1100);
 assign sub_590_52_n_31 = ~(n_1024 | n_1320);
 assign sub_590_52_n_29 = ~n_1349;
 assign sub_590_52_n_28 = ~{in1[0]};
 assign sub_590_52_n_23 = ~(sub_590_52_n_70 & ~sub_590_52_n_90);
 assign sub_590_52_n_22 = ~(sub_590_52_n_85 | (~sub_590_52_n_26 & sub_590_52_n_77));
 assign sub_590_52_n_21 = ~(sub_590_52_n_74 & ~sub_590_52_n_25);
 assign sub_590_52_n_20 = ~(sub_590_52_n_71 | (~sub_590_52_n_72 & sub_590_52_n_59));
 assign T_19_5_ = ~(sub_590_52_n_92 ^ sub_590_52_n_12);
 assign T_19_4_ = (sub_590_52_n_26 ^ sub_590_52_n_13);
 assign sub_590_52_n_17 = ~(sub_590_52_n_59 & ~sub_590_52_n_63);
 assign sub_590_52_n_16 = ~(sub_590_52_n_38 | ~sub_590_52_n_50);
 assign sub_590_52_n_15 = ~(sub_590_52_n_36 | ~sub_590_52_n_2);
 assign sub_590_52_n_14 = ~(sub_590_52_n_7 & ~sub_590_52_n_46);
 assign sub_590_52_n_13 = ~(sub_590_52_n_1 & ~sub_590_52_n_45);
 assign sub_590_52_n_12 = ~(sub_590_52_n_3 & ~sub_590_52_n_44);
 assign sub_590_52_n_11 = ~(sub_590_52_n_24 | ~sub_590_52_n_8);
 assign sub_590_52_n_10 = ~(sub_590_52_n_49 | ~sub_590_52_n_42);
 assign sub_590_52_n_9 = ~(sub_590_52_n_37 | ~sub_590_52_n_41);
 assign sub_590_52_n_8 = ~(R_20_9_ & ~n_1344);
 assign sub_590_52_n_7 = ~(R_20_7_ & ~n_1216);
 assign sub_590_52_n_6 = ~(R_20_6_ & ~n_1166);
 assign sub_590_52_n_5 = ~(R_20_1_ & ~n_1100);
 assign sub_590_52_n_4 = ~(n_1095 & ~R_20_5_);
 assign sub_590_52_n_3 = ~(R_20_4_ & ~n_1048);
 assign sub_590_52_n_2 = ~(R_20_8_ & ~n_1161);
 assign sub_590_52_n_1 = ~(R_20_3_ & ~n_1339);
 assign sub_590_52_n_0 = (R_20_0_ | sub_590_52_n_29);
 assign T_18_13_ = ((sub_620_51_n_115 & sub_620_51_n_19) | ~(sub_620_51_n_115 | sub_620_51_n_19));
 assign T_18_11_ = ~((sub_620_51_n_111 | sub_620_51_n_11) & ~(sub_620_51_n_111 & sub_620_51_n_11));
 assign sub_620_51_n_115 = ~(sub_620_51_n_48 | (~sub_620_51_n_41 & sub_620_51_n_108));
 assign T_18_12_ = ~((sub_620_51_n_108 | sub_620_51_n_12) & ~(sub_620_51_n_108 & sub_620_51_n_12));
 assign T_18_7_ = ((sub_620_51_n_106 & sub_620_51_n_14) | ~(sub_620_51_n_106 | sub_620_51_n_14));
 assign T_18_32_ = ~(sub_620_51_n_107 & ~sub_620_51_n_93);
 assign sub_620_51_n_111 = ~(sub_620_51_n_0 & (~sub_620_51_n_51 | sub_620_51_n_23));
 assign T_18_10_ = ~((sub_620_51_n_23 | sub_620_51_n_10) & ~(sub_620_51_n_23 & sub_620_51_n_10));
 assign T_18_9_ = ~((sub_620_51_n_16 | sub_620_51_n_13) & ~(sub_620_51_n_16 & sub_620_51_n_13));
 assign sub_620_51_n_108 = ~(sub_620_51_n_103 & ~sub_620_51_n_85);
 assign sub_620_51_n_107 = ~(sub_620_51_n_103 & ~sub_620_51_n_94);
 assign sub_620_51_n_106 = ~(sub_620_51_n_49 | (sub_620_51_n_22 & n_990));
 assign T_18_6_ = ((sub_620_51_n_22 & sub_620_51_n_67) | ~(sub_620_51_n_22 | sub_620_51_n_67));
 assign T_18_5_ = ((sub_620_51_n_100 & sub_620_51_n_65) | ~(sub_620_51_n_100 | sub_620_51_n_65));
 assign sub_620_51_n_103 = ~(sub_620_51_n_101 & ~sub_620_51_n_70);
 assign T_18_8_ = ((sub_620_51_n_98 & sub_620_51_n_15) | ~(sub_620_51_n_98 | sub_620_51_n_15));
 assign sub_620_51_n_101 = ~(sub_620_51_n_98 | ~sub_620_51_n_66);
 assign sub_620_51_n_100 = ~(n_1012 | (~n_1006 & sub_620_51_n_97));
 assign T_18_3_ = ~((sub_620_51_n_96 | sub_620_51_n_71) & ~(sub_620_51_n_96 & sub_620_51_n_71));
 assign sub_620_51_n_98 = ~(sub_620_51_n_86 | (sub_620_51_n_92 & sub_620_51_n_81));
 assign sub_620_51_n_97 = ~(sub_620_51_n_75 & (sub_620_51_n_91 | sub_620_51_n_62));
 assign sub_620_51_n_96 = ~(sub_620_51_n_47 & (~n_1002 | sub_620_51_n_88));
 assign T_18_2_ = ((sub_620_51_n_89 & sub_620_51_n_63) | ~(sub_620_51_n_89 | sub_620_51_n_63));
 assign sub_620_51_n_94 = ~(sub_620_51_n_84 & sub_620_51_n_82);
 assign sub_620_51_n_93 = ~(sub_620_51_n_80 & sub_620_51_n_90);
 assign sub_620_51_n_92 = ~(sub_620_51_n_73 | (sub_620_51_n_83 & sub_620_51_n_64));
 assign sub_620_51_n_91 = ~(n_1011 & ~n_1007);
 assign sub_620_51_n_90 = ~(sub_620_51_n_82 & ~sub_620_51_n_79);
 assign sub_620_51_n_89 = ~sub_620_51_n_88;
 assign sub_620_51_n_88 = ~(sub_620_51_n_24 | ~n_1010);
 assign T_18_1_ = ((sub_620_51_n_72 & n_1128) | ~(sub_620_51_n_72 | n_1128));
 assign sub_620_51_n_86 = ~(sub_620_51_n_76 & (sub_620_51_n_17 | sub_620_51_n_68));
 assign sub_620_51_n_85 = ~sub_620_51_n_84;
 assign sub_620_51_n_84 = ~(sub_620_51_n_74 | (sub_620_51_n_78 & sub_620_51_n_69));
 assign sub_620_51_n_83 = ~n_1011;
 assign sub_620_51_n_30 = ~(sub_620_51_n_40 & ~n_1127);
 assign sub_620_51_n_82 = ~(sub_620_51_n_77 & ~sub_620_51_n_45);
 assign sub_620_51_n_81 = ~(sub_620_51_n_68 | (sub_620_51_n_64 & sub_620_51_n_62));
 assign sub_620_51_n_80 = (sub_620_51_n_56 & (sub_620_51_n_57 & (sub_620_51_n_55 & sub_620_51_n_58)));
 assign sub_620_51_n_79 = ~(sub_620_51_n_45 | (sub_620_51_n_41 | sub_620_51_n_26));
 assign sub_620_51_n_78 = ~(n_998 & (sub_620_51_n_2 | n_997));
 assign sub_620_51_n_77 = ~(sub_620_51_n_54 & (sub_620_51_n_4 | sub_620_51_n_26));
 assign sub_620_51_n_76 = ~(n_1014 | (sub_620_51_n_49 & n_1015));
 assign sub_620_51_n_75 = ~(sub_620_51_n_43 | (n_1001 & sub_620_51_n_38));
 assign sub_620_51_n_74 = ~(sub_620_51_n_3 & (sub_620_51_n_0 | sub_620_51_n_39));
 assign sub_620_51_n_73 = ~(sub_620_51_n_60 & sub_620_51_n_61);
 assign sub_620_51_n_70 = ~sub_620_51_n_69;
 assign sub_620_51_n_66 = ~(sub_620_51_n_29 | n_997);
 assign sub_620_51_n_72 = ~(n_1010 & n_1009);
 assign sub_620_51_n_71 = ~(n_1005 & sub_620_51_n_38);
 assign sub_620_51_n_69 = ~(sub_620_51_n_50 | sub_620_51_n_39);
 assign sub_620_51_n_68 = ~(n_990 & n_1015);
 assign sub_620_51_n_67 = ~(n_991 & n_990);
 assign sub_620_51_n_60 = ~(n_1007 & n_1005);
 assign T_18_0_ = ~(sub_620_51_n_36 & (~{in2[18]} | {in1[0]}));
 assign sub_620_51_n_58 = ~(n_1297 | (n_1361 | (n_830 | n_1273)));
 assign sub_620_51_n_57 = ~(n_1212 | (n_1366 | (n_1177 | n_1292)));
 assign sub_620_51_n_56 = ~(n_1136 | (n_1172 | (n_1031 | n_1302)));
 assign sub_620_51_n_55 = ~(n_1059 | (n_1371 | (n_1086 | n_1242)));
 assign sub_620_51_n_65 = ~(n_988 | n_993);
 assign sub_620_51_n_64 = ~(n_1001 | ~n_1005);
 assign sub_620_51_n_63 = ~(sub_620_51_n_47 & n_1002);
 assign sub_620_51_n_62 = ~(n_1009 & n_1002);
 assign sub_620_51_n_61 = ~(n_1006 | n_993);
 assign sub_620_51_n_51 = ~sub_620_51_n_50;
 assign sub_620_51_n_49 = ~n_991;
 assign sub_620_51_n_48 = ~sub_620_51_n_4;
 assign sub_620_51_n_47 = ~n_1001;
 assign sub_620_51_n_54 = ~(n_995 & ~n_1259);
 assign sub_620_51_n_53 = ~(R_19_3_ | ~n_1339);
 assign sub_620_51_n_52 = ~(R_19_4_ | ~n_1048);
 assign sub_620_51_n_50 = ~(n_1016 | ~n_1345);
 assign sub_620_51_n_29 = ~(n_999 | ~n_1217);
 assign sub_620_51_n_28 = ~(sub_620_51_n_33 & R_19_5_);
 assign sub_620_51_n_46 = ~(n_1100 | sub_620_51_n_35);
 assign sub_620_51_n_43 = ~n_1005;
 assign sub_620_51_n_38 = ~n_1007;
 assign sub_620_51_n_45 = (n_1182 | n_1091);
 assign sub_620_51_n_44 = ~(R_19_8_ & ~n_1161);
 assign sub_620_51_n_42 = ~(R_19_8_ | ~n_1161);
 assign sub_620_51_n_41 = ~(n_992 | ~n_1026);
 assign sub_620_51_n_40 = ~(R_19_0_ & ~n_1349);
 assign sub_620_51_n_39 = ~(n_994 | ~n_1065);
 assign sub_620_51_n_37 = ~(R_19_2_ | ~n_1112);
 assign sub_620_51_n_36 = ~({in1[0]} & ~{in2[18]});
 assign sub_620_51_n_35 = ~R_19_1_;
 assign sub_620_51_n_34 = ~n_1166;
 assign sub_620_51_n_33 = ~n_1095;
 assign sub_620_51_n_32 = ~n_1112;
 assign sub_620_51_n_26 = ~(n_995 | ~n_1259);
 assign sub_620_51_n_27 = ~(sub_620_51_n_32 & R_19_2_);
 assign sub_620_51_n_25 = (sub_620_51_n_34 & R_19_6_);
 assign sub_620_51_n_24 = (n_1128 & n_1009);
 assign sub_620_51_n_23 = ~(sub_620_51_n_101 | sub_620_51_n_78);
 assign sub_620_51_n_22 = ~(sub_620_51_n_20 & sub_620_51_n_17);
 assign T_18_4_ = ~(sub_620_51_n_97 ^ sub_620_51_n_18);
 assign sub_620_51_n_20 = ~(sub_620_51_n_97 & sub_620_51_n_61);
 assign sub_620_51_n_19 = ~(sub_620_51_n_26 | ~sub_620_51_n_54);
 assign sub_620_51_n_18 = (n_1012 | n_1006);
 assign sub_620_51_n_17 = ~(n_988 | (~n_993 & n_1012));
 assign sub_620_51_n_16 = ~(sub_620_51_n_2 & (sub_620_51_n_29 | sub_620_51_n_98));
 assign sub_620_51_n_15 = ~(sub_620_51_n_29 | ~sub_620_51_n_2);
 assign sub_620_51_n_14 = ~(n_1014 | ~n_1015);
 assign sub_620_51_n_13 = ~(n_998 & ~n_997);
 assign sub_620_51_n_12 = ~(sub_620_51_n_4 & ~sub_620_51_n_41);
 assign sub_620_51_n_11 = ~(sub_620_51_n_3 & ~sub_620_51_n_39);
 assign sub_620_51_n_10 = ~(sub_620_51_n_50 | ~sub_620_51_n_0);
 assign sub_620_51_n_9 = ~(n_1048 | ~R_19_4_);
 assign sub_620_51_n_8 = ~(n_1349 & ~R_19_0_);
 assign sub_620_51_n_7 = (R_19_6_ | sub_620_51_n_34);
 assign sub_620_51_n_6 = ~(n_1339 | ~R_19_3_);
 assign sub_620_51_n_5 = ~(sub_620_51_n_35 & n_1100);
 assign sub_620_51_n_4 = ~(n_992 & ~n_1026);
 assign sub_620_51_n_3 = ~(n_994 & ~n_1065);
 assign sub_620_51_n_2 = ~(n_999 & ~n_1217);
 assign sub_620_51_n_1 = (R_19_5_ | sub_620_51_n_33);
 assign sub_620_51_n_0 = ~(n_1016 & ~n_1345);
 assign T_17_14_ = ~((sub_650_50_n_27 | sub_650_50_n_17) & ~(sub_650_50_n_27 & sub_650_50_n_17));
 assign T_17_13_ = ((sub_650_50_n_74 & ~sub_650_50_n_126) | (sub_650_50_n_23 & sub_650_50_n_126));
 assign T_17_11_ = ((sub_650_50_n_31 & sub_650_50_n_18) | ~(sub_650_50_n_31 | sub_650_50_n_18));
 assign sub_650_50_n_126 = ~(sub_650_50_n_53 & (~sub_650_50_n_3 | sub_650_50_n_119));
 assign T_17_12_ = ((sub_650_50_n_118 & sub_650_50_n_67) | ~(sub_650_50_n_118 | sub_650_50_n_67));
 assign T_17_10_ = ((sub_650_50_n_117 & sub_650_50_n_75) | ~(sub_650_50_n_117 | sub_650_50_n_75));
 assign T_17_9_ = ((sub_650_50_n_116 & sub_650_50_n_78) | ~(sub_650_50_n_116 | sub_650_50_n_78));
 assign T_17_7_ = ~((sub_650_50_n_15 | sub_650_50_n_13) & ~(sub_650_50_n_15 & sub_650_50_n_13));
 assign T_17_32_ = ~(sub_650_50_n_120 & ~sub_650_50_n_90);
 assign sub_650_50_n_120 = ~((sub_650_50_n_104 & sub_650_50_n_26) | (sub_650_50_n_111 & sub_650_50_n_103));
 assign sub_650_50_n_118 = ~sub_650_50_n_119;
 assign sub_650_50_n_119 = ~(sub_650_50_n_95 | (~sub_650_50_n_88 & sub_650_50_n_30));
 assign sub_650_50_n_117 = ~(sub_650_50_n_28 & (sub_650_50_n_98 | (sub_650_50_n_108 & sub_650_50_n_92)));
 assign sub_650_50_n_116 = ~(sub_650_50_n_55 & (~sub_650_50_n_57 | sub_650_50_n_110));
 assign T_17_8_ = ((sub_650_50_n_30 & sub_650_50_n_70) | ~(sub_650_50_n_30 | sub_650_50_n_70));
 assign T_17_6_ = ((sub_650_50_n_112 & sub_650_50_n_21) | ~(sub_650_50_n_112 | sub_650_50_n_21));
 assign T_17_3_ = ~((sub_650_50_n_12 | sub_650_50_n_16) & ~(sub_650_50_n_12 & sub_650_50_n_16));
 assign sub_650_50_n_112 = ~(sub_650_50_n_107 | ~sub_650_50_n_84);
 assign sub_650_50_n_111 = ~(sub_650_50_n_106 | sub_650_50_n_99);
 assign sub_650_50_n_110 = ~sub_650_50_n_30;
 assign T_17_4_ = ((sub_650_50_n_101 & sub_650_50_n_20) | ~(sub_650_50_n_101 | sub_650_50_n_20));
 assign sub_650_50_n_108 = ~sub_650_50_n_107;
 assign sub_650_50_n_107 = ~(sub_650_50_n_101 | ~sub_650_50_n_68);
 assign sub_650_50_n_106 = ~(sub_650_50_n_101 | sub_650_50_n_87);
 assign T_17_2_ = ~((sub_650_50_n_97 | sub_650_50_n_24) & ~(sub_650_50_n_97 & sub_650_50_n_24));
 assign sub_650_50_n_104 = ~(sub_650_50_n_29 & (~sub_650_50_n_88 | sub_650_50_n_95));
 assign sub_650_50_n_103 = ~(sub_650_50_n_95 | sub_650_50_n_94);
 assign sub_650_50_n_102 = ~(sub_650_50_n_97 & ~sub_650_50_n_59);
 assign sub_650_50_n_101 = ~(sub_650_50_n_79 | (sub_650_50_n_81 & sub_650_50_n_91));
 assign sub_650_50_n_100 = ~(sub_650_50_n_82 | (sub_650_50_n_83 & sub_650_50_n_37));
 assign sub_650_50_n_99 = ~(sub_650_50_n_93 & (sub_650_50_n_84 | sub_650_50_n_66));
 assign sub_650_50_n_98 = ~(sub_650_50_n_76 & (sub_650_50_n_82 | sub_650_50_n_37));
 assign sub_650_50_n_97 = ~(sub_650_50_n_4 & (sub_650_50_n_49 | sub_650_50_n_50));
 assign T_17_1_ = ((sub_650_50_n_19 & sub_650_50_n_89) | ~(sub_650_50_n_19 | sub_650_50_n_89));
 assign sub_650_50_n_95 = ~(sub_650_50_n_86 | (sub_650_50_n_80 & sub_650_50_n_73));
 assign sub_650_50_n_94 = ~(sub_650_50_n_85 | ~sub_650_50_n_77);
 assign sub_650_50_n_93 = ~(sub_650_50_n_82 | sub_650_50_n_71);
 assign sub_650_50_n_92 = ~(sub_650_50_n_83 | sub_650_50_n_82);
 assign sub_650_50_n_91 = ~(sub_650_50_n_49 & sub_650_50_n_4);
 assign sub_650_50_n_90 = ~(sub_650_50_n_60 & (sub_650_50_n_65 & (sub_650_50_n_61 & sub_650_50_n_62)));
 assign sub_650_50_n_89 = ~sub_650_50_n_49;
 assign sub_650_50_n_87 = ~(sub_650_50_n_68 & sub_650_50_n_37);
 assign sub_650_50_n_86 = ~(sub_650_50_n_69 | ~sub_650_50_n_45);
 assign sub_650_50_n_88 = ~(sub_650_50_n_76 & sub_650_50_n_69);
 assign sub_650_50_n_83 = ~sub_650_50_n_84;
 assign sub_650_50_n_81 = ~(sub_650_50_n_48 | (sub_650_50_n_32 | sub_650_50_n_50));
 assign sub_650_50_n_80 = ~(sub_650_50_n_6 | ~sub_650_50_n_58);
 assign sub_650_50_n_79 = ~(sub_650_50_n_7 & (sub_650_50_n_33 | sub_650_50_n_32));
 assign sub_650_50_n_85 = ~(sub_650_50_n_10 | (~sub_650_50_n_54 & sub_650_50_n_2));
 assign sub_650_50_n_84 = ~(sub_650_50_n_64 | ~sub_650_50_n_9);
 assign sub_650_50_n_82 = ~(sub_650_50_n_5 & (sub_650_50_n_8 | sub_650_50_n_41));
 assign sub_650_50_n_74 = ~sub_650_50_n_23;
 assign sub_650_50_n_78 = ~(sub_650_50_n_0 & sub_650_50_n_52);
 assign sub_650_50_n_77 = ~(sub_650_50_n_46 | ~sub_650_50_n_39);
 assign sub_650_50_n_76 = ~(sub_650_50_n_56 | sub_650_50_n_51);
 assign sub_650_50_n_75 = ~(sub_650_50_n_58 & sub_650_50_n_44);
 assign sub_650_50_n_73 = ~(sub_650_50_n_11 & sub_650_50_n_52);
 assign sub_650_50_n_72 = ~(sub_650_50_n_3 & ~sub_650_50_n_54);
 assign sub_650_50_n_71 = ~(sub_650_50_n_1 | ~sub_650_50_n_39);
 assign sub_650_50_n_66 = ~sub_650_50_n_37;
 assign sub_650_50_n_65 = ~(n_1212 | (n_1366 | (n_1177 | n_1292)));
 assign sub_650_50_n_64 = ~(sub_650_50_n_35 | sub_650_50_n_42);
 assign T_17_0_ = (sub_650_50_n_49 | (n_1319 & n_1056));
 assign sub_650_50_n_62 = ~(n_1297 | (n_1361 | (n_830 | n_1273)));
 assign sub_650_50_n_61 = ~(n_1059 | (n_1371 | (n_1086 | n_1242)));
 assign sub_650_50_n_60 = ~(n_1136 | (n_1172 | (n_1031 | n_1302)));
 assign sub_650_50_n_70 = ~(sub_650_50_n_55 & sub_650_50_n_57);
 assign sub_650_50_n_69 = ~(sub_650_50_n_43 | sub_650_50_n_47);
 assign sub_650_50_n_68 = ~(sub_650_50_n_36 | sub_650_50_n_42);
 assign sub_650_50_n_67 = ~(sub_650_50_n_53 & sub_650_50_n_3);
 assign sub_650_50_n_37 = ~(sub_650_50_n_34 | sub_650_50_n_41);
 assign sub_650_50_n_57 = ~sub_650_50_n_56;
 assign sub_650_50_n_55 = ~sub_650_50_n_11;
 assign sub_650_50_n_53 = ~sub_650_50_n_2;
 assign sub_650_50_n_52 = ~sub_650_50_n_51;
 assign sub_650_50_n_48 = ~(R_18_1_ | ~n_1101);
 assign sub_650_50_n_59 = ~(R_18_1_ | ~n_1101);
 assign sub_650_50_n_36 = ~(R_18_3_ | ~n_1340);
 assign sub_650_50_n_58 = ~(R_18_9_ & ~n_1345);
 assign sub_650_50_n_56 = ~(R_18_7_ | ~n_1217);
 assign sub_650_50_n_35 = ~(R_18_3_ & ~n_1340);
 assign sub_650_50_n_54 = ~(R_18_12_ | ~n_1259);
 assign sub_650_50_n_51 = ~(R_18_8_ | ~n_1162);
 assign sub_650_50_n_50 = ~(R_18_0_ | ~n_1350);
 assign sub_650_50_n_49 = ~(n_1056 | n_1319);
 assign sub_650_50_n_44 = ~sub_650_50_n_43;
 assign sub_650_50_n_47 = ~(R_18_10_ | ~n_1065);
 assign sub_650_50_n_46 = ~(R_18_13_ | ~n_1182);
 assign sub_650_50_n_45 = ~(R_18_10_ & ~n_1065);
 assign sub_650_50_n_34 = ~(R_18_5_ | ~n_1096);
 assign sub_650_50_n_43 = ~(R_18_9_ | ~n_1345);
 assign sub_650_50_n_42 = ~(R_18_4_ | ~n_1049);
 assign sub_650_50_n_41 = ~(R_18_6_ | ~n_1167);
 assign sub_650_50_n_33 = ~(R_18_1_ & ~n_1101);
 assign sub_650_50_n_40 = ~{in1[0]};
 assign sub_650_50_n_39 = ~n_1091;
 assign sub_650_50_n_32 = ~(R_18_2_ | ~n_1113);
 assign sub_650_50_n_31 = ~(sub_650_50_n_58 & ~(sub_650_50_n_44 & sub_650_50_n_117));
 assign sub_650_50_n_30 = ~(sub_650_50_n_100 & ~sub_650_50_n_106);
 assign sub_650_50_n_29 = ~(sub_650_50_n_72 | ~sub_650_50_n_77);
 assign sub_650_50_n_28 = (sub_650_50_n_73 & sub_650_50_n_0);
 assign sub_650_50_n_27 = ~(sub_650_50_n_85 & (sub_650_50_n_72 | sub_650_50_n_119));
 assign sub_650_50_n_26 = ~(sub_650_50_n_94 | sub_650_50_n_71);
 assign T_17_5_ = ~(sub_650_50_n_22 ^ sub_650_50_n_14);
 assign sub_650_50_n_24 = ~(sub_650_50_n_33 & ~sub_650_50_n_59);
 assign sub_650_50_n_23 = (sub_650_50_n_10 | sub_650_50_n_54);
 assign sub_650_50_n_22 = ~(sub_650_50_n_35 & (sub_650_50_n_36 | sub_650_50_n_101));
 assign sub_650_50_n_21 = ~(sub_650_50_n_34 | ~sub_650_50_n_8);
 assign sub_650_50_n_20 = ~(sub_650_50_n_36 | ~sub_650_50_n_35);
 assign sub_650_50_n_19 = ~(sub_650_50_n_4 & ~sub_650_50_n_50);
 assign sub_650_50_n_18 = ~(sub_650_50_n_45 & ~sub_650_50_n_47);
 assign sub_650_50_n_17 = ~(sub_650_50_n_1 & ~sub_650_50_n_46);
 assign sub_650_50_n_16 = ~(sub_650_50_n_7 & ~sub_650_50_n_32);
 assign sub_650_50_n_15 = ~(sub_650_50_n_8 & (sub_650_50_n_34 | sub_650_50_n_112));
 assign sub_650_50_n_14 = ~(sub_650_50_n_9 & ~sub_650_50_n_42);
 assign sub_650_50_n_13 = ~(sub_650_50_n_5 & ~sub_650_50_n_41);
 assign sub_650_50_n_12 = ~(sub_650_50_n_102 & sub_650_50_n_33);
 assign sub_650_50_n_11 = ~(n_1217 | ~R_18_7_);
 assign sub_650_50_n_10 = ~(n_1259 | ~R_18_12_);
 assign sub_650_50_n_9 = ~(R_18_4_ & ~n_1049);
 assign sub_650_50_n_8 = ~(R_18_5_ & ~n_1096);
 assign sub_650_50_n_7 = ~(R_18_2_ & ~n_1113);
 assign sub_650_50_n_6 = ~(sub_650_50_n_0 & (~R_18_10_ | n_1065));
 assign sub_650_50_n_5 = ~(R_18_6_ & ~n_1167);
 assign sub_650_50_n_4 = ~(R_18_0_ & ~n_1350);
 assign sub_650_50_n_3 = ~(n_1026 & ~R_18_11_);
 assign sub_650_50_n_2 = ~(n_1026 | ~R_18_11_);
 assign sub_650_50_n_1 = ~(R_18_13_ & ~n_1182);
 assign sub_650_50_n_0 = ~(R_18_8_ & ~n_1162);
 assign T_16_15_ = ((sub_680_49_n_19 & sub_680_49_n_12) | ~(sub_680_49_n_19 | sub_680_49_n_12));
 assign T_16_13_ = ((sub_680_49_n_144 & sub_680_49_n_10) | ~(sub_680_49_n_144 | sub_680_49_n_10));
 assign T_16_11_ = ((sub_680_49_n_143 & sub_680_49_n_14) | ~(sub_680_49_n_143 | sub_680_49_n_14));
 assign sub_680_49_n_144 = ~(sub_680_49_n_56 & (~sub_680_49_n_42 | sub_680_49_n_133));
 assign sub_680_49_n_143 = ~(sub_680_49_n_1 & (~sub_680_49_n_59 | sub_680_49_n_17));
 assign T_16_14_ = ((sub_680_49_n_135 & sub_680_49_n_86) | ~(sub_680_49_n_135 | sub_680_49_n_86));
 assign T_16_12_ = ((sub_680_49_n_134 & sub_680_49_n_87) | ~(sub_680_49_n_134 | sub_680_49_n_87));
 assign T_16_10_ = ((sub_680_49_n_25 & sub_680_49_n_84) | ~(sub_680_49_n_25 | sub_680_49_n_84));
 assign T_16_9_ = ((sub_680_49_n_132 & sub_680_49_n_13) | ~(sub_680_49_n_132 | sub_680_49_n_13));
 assign T_16_7_ = ~((sub_680_49_n_11 | sub_680_49_n_89) & ~(sub_680_49_n_11 & sub_680_49_n_89));
 assign T_16_32_ = ~(sub_680_49_n_136 & ~sub_680_49_n_102);
 assign sub_680_49_n_136 = ~(sub_680_49_n_113 & (sub_680_49_n_21 & sub_680_49_n_127));
 assign sub_680_49_n_135 = ~(sub_680_49_n_119 & (sub_680_49_n_125 | sub_680_49_n_18));
 assign sub_680_49_n_134 = ~sub_680_49_n_133;
 assign sub_680_49_n_133 = ~(sub_680_49_n_108 | (~sub_680_49_n_100 & sub_680_49_n_126));
 assign sub_680_49_n_25 = ~sub_680_49_n_17;
 assign sub_680_49_n_132 = ~(sub_680_49_n_5 & (~sub_680_49_n_44 | sub_680_49_n_125));
 assign T_16_6_ = ~((sub_680_49_n_124 | sub_680_49_n_88) & ~(sub_680_49_n_124 & sub_680_49_n_88));
 assign T_16_5_ = ~((sub_680_49_n_123 | sub_680_49_n_85) & ~(sub_680_49_n_123 & sub_680_49_n_85));
 assign T_16_8_ = ~((sub_680_49_n_126 | sub_680_49_n_74) & ~(sub_680_49_n_126 & sub_680_49_n_74));
 assign sub_680_49_n_128 = ~(sub_680_49_n_124 & ~sub_680_49_n_38);
 assign sub_680_49_n_127 = ~(sub_680_49_n_126 & sub_680_49_n_16);
 assign sub_680_49_n_125 = ~sub_680_49_n_126;
 assign sub_680_49_n_126 = ~(sub_680_49_n_121 & sub_680_49_n_110);
 assign sub_680_49_n_124 = ~(sub_680_49_n_120 & ~sub_680_49_n_95);
 assign sub_680_49_n_123 = ~(sub_680_49_n_48 & (~sub_680_49_n_50 | sub_680_49_n_117));
 assign T_16_4_ = ~((sub_680_49_n_118 | sub_680_49_n_75) & ~(sub_680_49_n_118 & sub_680_49_n_75));
 assign sub_680_49_n_121 = ~(sub_680_49_n_112 & (sub_680_49_n_90 & sub_680_49_n_103));
 assign sub_680_49_n_120 = ~(sub_680_49_n_116 & ~sub_680_49_n_69);
 assign sub_680_49_n_119 = ~(sub_680_49_n_94 | (sub_680_49_n_108 & sub_680_49_n_82));
 assign sub_680_49_n_118 = ~sub_680_49_n_117;
 assign sub_680_49_n_117 = ~sub_680_49_n_116;
 assign sub_680_49_n_116 = ~(sub_680_49_n_91 & (sub_680_49_n_111 | sub_680_49_n_72));
 assign sub_680_49_n_115 = ~(sub_680_49_n_7 & (~sub_680_49_n_37 | sub_680_49_n_111));
 assign T_16_2_ = ~((sub_680_49_n_111 | sub_680_49_n_83) & ~(sub_680_49_n_111 & sub_680_49_n_83));
 assign sub_680_49_n_113 = ~(sub_680_49_n_82 & (sub_680_49_n_79 & sub_680_49_n_108));
 assign sub_680_49_n_112 = ~(sub_680_49_n_105 & (sub_680_49_n_7 & sub_680_49_n_20));
 assign sub_680_49_n_111 = ~(sub_680_49_n_106 | ~sub_680_49_n_60);
 assign sub_680_49_n_110 = ~(sub_680_49_n_96 | (sub_680_49_n_95 & sub_680_49_n_68));
 assign T_16_1_ = ((sub_680_49_n_77 & n_1257) | ~(sub_680_49_n_77 | n_1257));
 assign sub_680_49_n_108 = ~(sub_680_49_n_107 & ~sub_680_49_n_93);
 assign sub_680_49_n_107 = ~(sub_680_49_n_101 & sub_680_49_n_81);
 assign sub_680_49_n_106 = ~sub_680_49_n_105;
 assign sub_680_49_n_105 = ~(n_1257 & sub_680_49_n_62);
 assign sub_680_49_n_104 = ~(sub_680_49_n_94 & sub_680_49_n_79);
 assign sub_680_49_n_103 = ~(sub_680_49_n_92 | sub_680_49_n_78);
 assign sub_680_49_n_102 = ~(sub_680_49_n_73 & (sub_680_49_n_70 & (sub_680_49_n_71 & sub_680_49_n_67)));
 assign sub_680_49_n_99 = ~(sub_680_49_n_2 & (sub_680_49_n_45 | sub_680_49_n_55));
 assign sub_680_49_n_98 = ~(sub_680_49_n_80 & sub_680_49_n_42);
 assign sub_680_49_n_97 = ~(sub_680_49_n_81 & ~sub_680_49_n_40);
 assign sub_680_49_n_96 = ~(sub_680_49_n_63 & (sub_680_49_n_23 | sub_680_49_n_39));
 assign sub_680_49_n_101 = ~(sub_680_49_n_8 & (sub_680_49_n_5 | sub_680_49_n_57));
 assign sub_680_49_n_100 = ~(sub_680_49_n_80 & sub_680_49_n_81);
 assign sub_680_49_n_93 = ~(sub_680_49_n_0 & (sub_680_49_n_1 | sub_680_49_n_61));
 assign sub_680_49_n_92 = ~(sub_680_49_n_64 | ~sub_680_49_n_7);
 assign sub_680_49_n_91 = ~(sub_680_49_n_36 | (sub_680_49_n_35 & sub_680_49_n_54));
 assign sub_680_49_n_90 = ~(sub_680_49_n_65 | (sub_680_49_n_53 & sub_680_49_n_9));
 assign sub_680_49_n_95 = ~(sub_680_49_n_3 & (sub_680_49_n_52 | sub_680_49_n_48));
 assign sub_680_49_n_94 = ~(sub_680_49_n_49 & (sub_680_49_n_56 | sub_680_49_n_40));
 assign sub_680_49_n_78 = ~(sub_680_49_n_24 & sub_680_49_n_6);
 assign sub_680_49_n_89 = ~(sub_680_49_n_63 & sub_680_49_n_4);
 assign sub_680_49_n_88 = ~(sub_680_49_n_23 & sub_680_49_n_6);
 assign sub_680_49_n_87 = ~(sub_680_49_n_56 & sub_680_49_n_42);
 assign sub_680_49_n_86 = ~(sub_680_49_n_45 & sub_680_49_n_47);
 assign sub_680_49_n_85 = ~(sub_680_49_n_3 & sub_680_49_n_24);
 assign sub_680_49_n_84 = ~(sub_680_49_n_1 & sub_680_49_n_59);
 assign sub_680_49_n_83 = ~(sub_680_49_n_35 | sub_680_49_n_22);
 assign sub_680_49_n_82 = ~(sub_680_49_n_41 | sub_680_49_n_40);
 assign sub_680_49_n_81 = ~(sub_680_49_n_58 | sub_680_49_n_61);
 assign sub_680_49_n_80 = ~(sub_680_49_n_43 | sub_680_49_n_57);
 assign sub_680_49_n_79 = ~(sub_680_49_n_46 | sub_680_49_n_55);
 assign sub_680_49_n_73 = ~(n_1136 | (n_1172 | (n_1031 | n_1302)));
 assign sub_680_49_n_72 = ~(sub_680_49_n_37 & sub_680_49_n_54);
 assign sub_680_49_n_71 = ~(n_1059 | (n_1371 | (n_1086 | n_1242)));
 assign sub_680_49_n_70 = ~(n_1212 | (n_1366 | (n_1177 | n_1292)));
 assign sub_680_49_n_69 = ~(sub_680_49_n_50 & sub_680_49_n_24);
 assign sub_680_49_n_68 = ~(sub_680_49_n_38 | sub_680_49_n_39);
 assign sub_680_49_n_67 = ~(n_1297 | (n_1361 | (n_830 | n_1273)));
 assign T_16_0_ = ~(sub_680_49_n_51 & (~{in2[16]} | {in1[0]}));
 assign sub_680_49_n_65 = ~(sub_680_49_n_50 & sub_680_49_n_4);
 assign sub_680_49_n_64 = ~(sub_680_49_n_22 & sub_680_49_n_9);
 assign sub_680_49_n_77 = ~(sub_680_49_n_60 & sub_680_49_n_62);
 assign sub_680_49_n_76 = ~(sub_680_49_n_9 & sub_680_49_n_54);
 assign sub_680_49_n_75 = ~(sub_680_49_n_48 & sub_680_49_n_50);
 assign sub_680_49_n_74 = ~(sub_680_49_n_5 & sub_680_49_n_44);
 assign sub_680_49_n_59 = ~sub_680_49_n_58;
 assign sub_680_49_n_54 = ~sub_680_49_n_53;
 assign sub_680_49_n_52 = ~sub_680_49_n_24;
 assign sub_680_49_n_63 = ~(sub_680_49_n_29 & R_17_6_);
 assign sub_680_49_n_62 = ~(sub_680_49_n_33 & ~sub_680_49_n_30);
 assign sub_680_49_n_61 = ~(R_17_10_ | ~n_1065);
 assign sub_680_49_n_60 = ~(sub_680_49_n_30 & R_17_0_);
 assign sub_680_49_n_58 = ~(R_17_9_ | ~n_1345);
 assign sub_680_49_n_57 = ~(R_17_8_ | ~n_1162);
 assign sub_680_49_n_56 = ~(R_17_11_ & ~n_1026);
 assign sub_680_49_n_55 = ~(R_17_14_ | ~n_1091);
 assign sub_680_49_n_53 = ~(R_17_2_ | ~n_1113);
 assign sub_680_49_n_24 = ~(sub_680_49_n_31 & ~sub_680_49_n_34);
 assign sub_680_49_n_51 = ~({in1[0]} & ~{in2[16]});
 assign sub_680_49_n_50 = ~(sub_680_49_n_27 & ~sub_680_49_n_32);
 assign sub_680_49_n_47 = ~sub_680_49_n_46;
 assign sub_680_49_n_44 = ~sub_680_49_n_43;
 assign sub_680_49_n_42 = ~sub_680_49_n_41;
 assign sub_680_49_n_39 = ~sub_680_49_n_4;
 assign sub_680_49_n_38 = ~sub_680_49_n_6;
 assign sub_680_49_n_37 = ~sub_680_49_n_22;
 assign sub_680_49_n_36 = ~sub_680_49_n_9;
 assign sub_680_49_n_35 = ~sub_680_49_n_7;
 assign sub_680_49_n_49 = ~(R_17_12_ & ~n_1259);
 assign sub_680_49_n_23 = ~(R_17_5_ & ~n_1096);
 assign sub_680_49_n_48 = ~(sub_680_49_n_28 & ~n_1340);
 assign sub_680_49_n_46 = ~(R_17_13_ | ~n_1182);
 assign sub_680_49_n_45 = ~(R_17_13_ & ~n_1182);
 assign sub_680_49_n_43 = ~(R_17_7_ | ~n_1217);
 assign sub_680_49_n_41 = ~(R_17_11_ | ~n_1026);
 assign sub_680_49_n_40 = ~(R_17_12_ | ~n_1259);
 assign sub_680_49_n_22 = ~(R_17_1_ | ~n_1101);
 assign sub_680_49_n_34 = ~n_1049;
 assign sub_680_49_n_33 = ~R_17_0_;
 assign sub_680_49_n_32 = ~n_1340;
 assign sub_680_49_n_31 = ~R_17_4_;
 assign sub_680_49_n_30 = ~n_1350;
 assign sub_680_49_n_29 = ~n_1167;
 assign sub_680_49_n_28 = ~sub_680_49_n_27;
 assign sub_680_49_n_27 = ~R_17_3_;
 assign sub_680_49_n_21 = ~(sub_680_49_n_99 | ~sub_680_49_n_104);
 assign sub_680_49_n_20 = (sub_680_49_n_60 & sub_680_49_n_9);
 assign sub_680_49_n_19 = ~(sub_680_49_n_45 & ~(sub_680_49_n_47 & sub_680_49_n_135));
 assign sub_680_49_n_18 = ~(sub_680_49_n_82 & ~sub_680_49_n_100);
 assign sub_680_49_n_17 = ~(sub_680_49_n_101 | (sub_680_49_n_80 & sub_680_49_n_126));
 assign sub_680_49_n_16 = ~(sub_680_49_n_98 | (sub_680_49_n_97 | ~sub_680_49_n_79));
 assign T_16_3_ = ~(sub_680_49_n_115 ^ sub_680_49_n_76);
 assign sub_680_49_n_14 = ~(sub_680_49_n_0 & ~sub_680_49_n_61);
 assign sub_680_49_n_13 = ~(sub_680_49_n_8 & ~sub_680_49_n_57);
 assign sub_680_49_n_12 = ~(sub_680_49_n_2 & ~sub_680_49_n_55);
 assign sub_680_49_n_11 = ~(sub_680_49_n_128 & sub_680_49_n_23);
 assign sub_680_49_n_10 = ~(sub_680_49_n_49 & ~sub_680_49_n_40);
 assign sub_680_49_n_9 = ~(R_17_2_ & ~n_1113);
 assign sub_680_49_n_8 = ~(R_17_8_ & ~n_1162);
 assign sub_680_49_n_7 = ~(R_17_1_ & ~n_1101);
 assign sub_680_49_n_6 = ~(n_1096 & ~R_17_5_);
 assign sub_680_49_n_5 = ~(R_17_7_ & ~n_1217);
 assign sub_680_49_n_4 = (R_17_6_ | sub_680_49_n_29);
 assign sub_680_49_n_3 = ~(sub_680_49_n_34 & ~sub_680_49_n_31);
 assign sub_680_49_n_2 = ~(R_17_14_ & ~n_1091);
 assign sub_680_49_n_1 = ~(R_17_9_ & ~n_1345);
 assign sub_680_49_n_0 = ~(R_17_10_ & ~n_1065);
 assign T_15_15_ = ~(sub_710_48_n_147 & sub_710_48_n_153);
 assign T_15_14_ = ((sub_710_48_n_148 & sub_710_48_n_92) | ~(sub_710_48_n_148 | sub_710_48_n_92));
 assign T_15_13_ = ((sub_710_48_n_21 & sub_710_48_n_91) | ~(sub_710_48_n_21 | sub_710_48_n_91));
 assign T_15_11_ = ((sub_710_48_n_146 & sub_710_48_n_87) | ~(sub_710_48_n_146 | sub_710_48_n_87));
 assign sub_710_48_n_153 = ~(sub_710_48_n_16 & ~sub_710_48_n_17);
 assign T_15_16_ = ~((sub_710_48_n_142 | sub_710_48_n_88) & ~(sub_710_48_n_142 & sub_710_48_n_88));
 assign T_15_7_ = ~((sub_710_48_n_137 | sub_710_48_n_14) & ~(sub_710_48_n_137 & sub_710_48_n_14));
 assign T_15_32_ = ~(sub_710_48_n_149 | ~sub_710_48_n_26);
 assign sub_710_48_n_149 = ~(sub_710_48_n_142 | ~sub_710_48_n_116);
 assign sub_710_48_n_148 = ~(sub_710_48_n_141 & ~sub_710_48_n_97);
 assign sub_710_48_n_147 = ~(sub_710_48_n_138 & ~sub_710_48_n_103);
 assign sub_710_48_n_146 = ~(sub_710_48_n_139 & ~sub_710_48_n_63);
 assign T_15_12_ = ~((sub_710_48_n_134 | sub_710_48_n_78) & ~(sub_710_48_n_134 & sub_710_48_n_78));
 assign T_15_10_ = ~((sub_710_48_n_132 | sub_710_48_n_20) & ~(sub_710_48_n_132 & sub_710_48_n_20));
 assign T_15_9_ = ((sub_710_48_n_29 & sub_710_48_n_89) | ~(sub_710_48_n_29 | sub_710_48_n_89));
 assign sub_710_48_n_142 = ~(sub_710_48_n_127 | (sub_710_48_n_117 | sub_710_48_n_121));
 assign sub_710_48_n_141 = ~(sub_710_48_n_134 & ~sub_710_48_n_85);
 assign sub_710_48_n_140 = ~(sub_710_48_n_134 & ~sub_710_48_n_46);
 assign sub_710_48_n_139 = ~(sub_710_48_n_132 & ~sub_710_48_n_66);
 assign sub_710_48_n_138 = ~(sub_710_48_n_133 & ~sub_710_48_n_25);
 assign sub_710_48_n_137 = ~(sub_710_48_n_1 & (~sub_710_48_n_6 | sub_710_48_n_24));
 assign T_15_6_ = ~((sub_710_48_n_128 | sub_710_48_n_90) & ~(sub_710_48_n_128 & sub_710_48_n_90));
 assign T_15_5_ = ((sub_710_48_n_126 & sub_710_48_n_93) | ~(sub_710_48_n_126 | sub_710_48_n_93));
 assign sub_710_48_n_134 = ~(sub_710_48_n_130 & ~sub_710_48_n_115);
 assign sub_710_48_n_133 = ~(sub_710_48_n_130 & ~sub_710_48_n_28);
 assign sub_710_48_n_132 = ~(sub_710_48_n_129 & ~sub_710_48_n_98);
 assign T_15_8_ = ((sub_710_48_n_123 & sub_710_48_n_75) | ~(sub_710_48_n_123 | sub_710_48_n_75));
 assign sub_710_48_n_130 = ~(sub_710_48_n_123 & ~sub_710_48_n_105);
 assign sub_710_48_n_129 = ~(sub_710_48_n_123 & ~sub_710_48_n_86);
 assign sub_710_48_n_128 = ~(sub_710_48_n_107 & (~sub_710_48_n_81 | sub_710_48_n_120));
 assign sub_710_48_n_127 = ~(sub_710_48_n_96 | (sub_710_48_n_105 | sub_710_48_n_122));
 assign sub_710_48_n_126 = ~(sub_710_48_n_65 & (~sub_710_48_n_57 | sub_710_48_n_120));
 assign T_15_4_ = ~((sub_710_48_n_34 | sub_710_48_n_80) & ~(sub_710_48_n_34 & sub_710_48_n_80));
 assign T_15_3_ = ((sub_710_48_n_119 & sub_710_48_n_18) | ~(sub_710_48_n_119 | sub_710_48_n_18));
 assign sub_710_48_n_123 = ~(sub_710_48_n_122 & sub_710_48_n_114);
 assign sub_710_48_n_122 = ~(sub_710_48_n_23 & (sub_710_48_n_95 & sub_710_48_n_108));
 assign sub_710_48_n_121 = ~(sub_710_48_n_113 & (sub_710_48_n_110 | sub_710_48_n_114));
 assign sub_710_48_n_120 = ~sub_710_48_n_34;
 assign sub_710_48_n_34 = ~(sub_710_48_n_30 & (~sub_710_48_n_73 | sub_710_48_n_27));
 assign sub_710_48_n_119 = ~(sub_710_48_n_62 & (sub_710_48_n_27 | sub_710_48_n_32));
 assign T_15_2_ = ~((sub_710_48_n_27 | sub_710_48_n_19) & ~(sub_710_48_n_27 & sub_710_48_n_19));
 assign sub_710_48_n_117 = ~((sub_710_48_n_96 | sub_710_48_n_99) & (sub_710_48_n_22 | sub_710_48_n_96));
 assign sub_710_48_n_116 = ~(sub_710_48_n_109 | sub_710_48_n_67);
 assign sub_710_48_n_115 = ~(sub_710_48_n_22 & sub_710_48_n_99);
 assign sub_710_48_n_114 = ~(sub_710_48_n_100 | (sub_710_48_n_106 & sub_710_48_n_15));
 assign sub_710_48_n_113 = ~(sub_710_48_n_102 | (sub_710_48_n_97 & sub_710_48_n_82));
 assign T_15_1_ = ~((sub_710_48_n_77 | n_1312) & ~(sub_710_48_n_77 & n_1312));
 assign sub_710_48_n_111 = ~(n_1312 & sub_710_48_n_9);
 assign sub_710_48_n_110 = ~(sub_710_48_n_104 & sub_710_48_n_94);
 assign sub_710_48_n_109 = ~(sub_710_48_n_72 & (sub_710_48_n_71 & (sub_710_48_n_74 & sub_710_48_n_69)));
 assign sub_710_48_n_108 = ~(sub_710_48_n_101 | sub_710_48_n_84);
 assign sub_710_48_n_107 = ~sub_710_48_n_106;
 assign sub_710_48_n_105 = ~sub_710_48_n_104;
 assign sub_710_48_n_103 = ~(sub_710_48_n_17 & sub_710_48_n_31);
 assign sub_710_48_n_102 = ~(sub_710_48_n_3 & (sub_710_48_n_31 | sub_710_48_n_43));
 assign sub_710_48_n_101 = ~(sub_710_48_n_79 | ~sub_710_48_n_32);
 assign sub_710_48_n_100 = ~(sub_710_48_n_2 & (sub_710_48_n_1 | sub_710_48_n_44));
 assign sub_710_48_n_106 = ~(sub_710_48_n_8 & (sub_710_48_n_65 | sub_710_48_n_58));
 assign sub_710_48_n_104 = ~(sub_710_48_n_86 | sub_710_48_n_76);
 assign sub_710_48_n_95 = ~(sub_710_48_n_56 | (sub_710_48_n_44 | (sub_710_48_n_60 & sub_710_48_n_55)));
 assign sub_710_48_n_99 = ~(sub_710_48_n_54 | (sub_710_48_n_63 & sub_710_48_n_7));
 assign sub_710_48_n_98 = ~(sub_710_48_n_10 & (sub_710_48_n_51 | sub_710_48_n_52));
 assign sub_710_48_n_97 = ~(sub_710_48_n_5 & (sub_710_48_n_64 | sub_710_48_n_50));
 assign sub_710_48_n_96 = ~(sub_710_48_n_83 & sub_710_48_n_70);
 assign sub_710_48_n_94 = ~(sub_710_48_n_46 | (sub_710_48_n_47 | sub_710_48_n_13));
 assign sub_710_48_n_84 = ~(sub_710_48_n_59 & sub_710_48_n_6);
 assign sub_710_48_n_83 = ~(sub_710_48_n_46 | sub_710_48_n_47);
 assign sub_710_48_n_82 = ~(sub_710_48_n_47 | sub_710_48_n_43);
 assign sub_710_48_n_93 = ~(sub_710_48_n_8 & sub_710_48_n_59);
 assign sub_710_48_n_92 = ~(sub_710_48_n_31 & sub_710_48_n_48);
 assign sub_710_48_n_91 = ~(sub_710_48_n_5 & sub_710_48_n_49);
 assign sub_710_48_n_90 = ~(sub_710_48_n_1 & sub_710_48_n_6);
 assign sub_710_48_n_89 = ~(sub_710_48_n_10 & sub_710_48_n_53);
 assign sub_710_48_n_88 = ~(sub_710_48_n_12 | sub_710_48_n_67);
 assign sub_710_48_n_87 = ~(sub_710_48_n_0 & sub_710_48_n_7);
 assign sub_710_48_n_86 = ~(sub_710_48_n_4 & sub_710_48_n_53);
 assign sub_710_48_n_85 = ~(sub_710_48_n_45 & ~sub_710_48_n_50);
 assign sub_710_48_n_74 = ~(n_1371 | (n_1086 | (n_1242 | n_1297)));
 assign sub_710_48_n_73 = ~(sub_710_48_n_32 | sub_710_48_n_60);
 assign sub_710_48_n_72 = ~(n_1172 | (n_1059 | (n_1031 | n_1302)));
 assign sub_710_48_n_71 = ~(n_1212 | (n_1366 | (n_1177 | n_1292)));
 assign sub_710_48_n_70 = ~(sub_710_48_n_50 | sub_710_48_n_43);
 assign sub_710_48_n_81 = ~(sub_710_48_n_56 | sub_710_48_n_58);
 assign sub_710_48_n_69 = ~(n_1361 | (n_830 | n_1273));
 assign T_15_0_ = ~(sub_710_48_n_61 & (~{in2[15]} | {in1[0]}));
 assign sub_710_48_n_80 = ~(sub_710_48_n_65 & sub_710_48_n_57);
 assign sub_710_48_n_79 = ~(sub_710_48_n_62 & sub_710_48_n_55);
 assign sub_710_48_n_78 = ~(sub_710_48_n_64 & sub_710_48_n_45);
 assign sub_710_48_n_77 = ~(sub_710_48_n_33 & sub_710_48_n_9);
 assign sub_710_48_n_76 = ~(sub_710_48_n_11 & sub_710_48_n_7);
 assign sub_710_48_n_75 = ~(sub_710_48_n_51 & sub_710_48_n_4);
 assign sub_710_48_n_66 = ~sub_710_48_n_11;
 assign sub_710_48_n_58 = ~sub_710_48_n_59;
 assign sub_710_48_n_57 = ~sub_710_48_n_56;
 assign sub_710_48_n_67 = ~(R_16_15_ | ~n_1136);
 assign sub_710_48_n_65 = ~(R_16_3_ & ~n_1340);
 assign sub_710_48_n_64 = ~(R_16_11_ & ~n_1026);
 assign sub_710_48_n_63 = ~(n_1345 | sub_710_48_n_41);
 assign sub_710_48_n_33 = ~(R_16_0_ & ~n_1350);
 assign sub_710_48_n_62 = ~(R_16_1_ & ~n_1101);
 assign sub_710_48_n_61 = ~({in1[0]} & ~{in2[15]});
 assign sub_710_48_n_60 = ~(R_16_2_ | ~n_1113);
 assign sub_710_48_n_59 = ~(sub_710_48_n_42 & ~sub_710_48_n_38);
 assign sub_710_48_n_56 = ~(R_16_3_ | ~n_1340);
 assign sub_710_48_n_55 = ~(R_16_2_ & ~n_1113);
 assign sub_710_48_n_54 = ~sub_710_48_n_0;
 assign sub_710_48_n_53 = ~sub_710_48_n_52;
 assign sub_710_48_n_49 = ~sub_710_48_n_50;
 assign sub_710_48_n_48 = ~sub_710_48_n_47;
 assign sub_710_48_n_45 = ~sub_710_48_n_46;
 assign sub_710_48_n_52 = ~(R_16_8_ | ~n_1162);
 assign sub_710_48_n_51 = ~(sub_710_48_n_39 & R_16_7_);
 assign sub_710_48_n_50 = ~(R_16_12_ | ~n_1259);
 assign sub_710_48_n_47 = ~(R_16_13_ | ~n_1182);
 assign sub_710_48_n_46 = ~(R_16_11_ | ~n_1026);
 assign sub_710_48_n_44 = ~(R_16_6_ | ~n_1167);
 assign sub_710_48_n_43 = ~(R_16_14_ | ~n_1091);
 assign sub_710_48_n_42 = ~R_16_4_;
 assign sub_710_48_n_41 = ~R_16_9_;
 assign sub_710_48_n_40 = ~n_1182;
 assign sub_710_48_n_39 = ~n_1217;
 assign sub_710_48_n_38 = ~n_1049;
 assign sub_710_48_n_37 = ~R_16_5_;
 assign sub_710_48_n_36 = ~R_16_10_;
 assign sub_710_48_n_32 = ~(R_16_1_ | ~n_1101);
 assign sub_710_48_n_31 = ~(sub_710_48_n_40 & R_16_13_);
 assign sub_710_48_n_30 = (sub_710_48_n_55 & (sub_710_48_n_62 | sub_710_48_n_60));
 assign sub_710_48_n_29 = ~(sub_710_48_n_51 & ~(sub_710_48_n_4 & sub_710_48_n_123));
 assign sub_710_48_n_28 = (sub_710_48_n_115 | sub_710_48_n_97);
 assign sub_710_48_n_27 = (sub_710_48_n_111 & sub_710_48_n_33);
 assign sub_710_48_n_26 = ~(sub_710_48_n_12 & ~sub_710_48_n_109);
 assign sub_710_48_n_25 = ~(sub_710_48_n_48 & (~sub_710_48_n_85 | sub_710_48_n_97));
 assign sub_710_48_n_24 = ~(sub_710_48_n_106 | (sub_710_48_n_81 & sub_710_48_n_34));
 assign sub_710_48_n_23 = ~(sub_710_48_n_111 & (sub_710_48_n_33 & ~sub_710_48_n_79));
 assign sub_710_48_n_22 = ~(sub_710_48_n_98 & ~sub_710_48_n_76);
 assign sub_710_48_n_21 = ~(sub_710_48_n_140 & sub_710_48_n_64);
 assign sub_710_48_n_20 = ~(sub_710_48_n_11 & ~sub_710_48_n_63);
 assign sub_710_48_n_19 = ~(sub_710_48_n_32 | ~sub_710_48_n_62);
 assign sub_710_48_n_18 = ~(sub_710_48_n_55 & ~sub_710_48_n_60);
 assign sub_710_48_n_17 = ~(sub_710_48_n_43 | ~sub_710_48_n_3);
 assign sub_710_48_n_16 = ~(sub_710_48_n_138 & sub_710_48_n_31);
 assign sub_710_48_n_15 = ~(sub_710_48_n_44 | ~sub_710_48_n_6);
 assign sub_710_48_n_14 = ~(sub_710_48_n_2 & ~sub_710_48_n_44);
 assign sub_710_48_n_13 = ~(sub_710_48_n_49 & ~sub_710_48_n_43);
 assign sub_710_48_n_12 = ~(n_1136 | ~R_16_15_);
 assign sub_710_48_n_11 = ~(sub_710_48_n_41 & n_1345);
 assign sub_710_48_n_10 = ~(R_16_8_ & ~n_1162);
 assign sub_710_48_n_9 = ~(n_1350 & ~R_16_0_);
 assign sub_710_48_n_8 = ~(sub_710_48_n_38 & ~sub_710_48_n_42);
 assign sub_710_48_n_7 = ~(sub_710_48_n_36 & n_1065);
 assign sub_710_48_n_6 = ~(sub_710_48_n_37 & n_1096);
 assign sub_710_48_n_5 = ~(R_16_12_ & ~n_1259);
 assign sub_710_48_n_4 = (R_16_7_ | sub_710_48_n_39);
 assign sub_710_48_n_3 = ~(R_16_14_ & ~n_1091);
 assign sub_710_48_n_2 = ~(R_16_6_ & ~n_1167);
 assign sub_710_48_n_1 = (sub_710_48_n_37 | n_1096);
 assign sub_710_48_n_0 = (sub_710_48_n_36 | n_1065);
 assign T_14_15_ = ((sub_740_47_n_143 & sub_740_47_n_22) | ~(sub_740_47_n_143 | sub_740_47_n_22));
 assign sub_740_47_n_143 = ~(sub_740_47_n_138 & ~sub_740_47_n_40);
 assign T_14_17_ = ~((sub_740_47_n_21 | sub_740_47_n_85) & ~(sub_740_47_n_21 & sub_740_47_n_85));
 assign T_14_14_ = ((sub_740_47_n_135 & sub_740_47_n_18) | ~(sub_740_47_n_135 | sub_740_47_n_18));
 assign T_14_13_ = ((sub_740_47_n_134 & sub_740_47_n_12) | ~(sub_740_47_n_134 | sub_740_47_n_12));
 assign T_14_11_ = ((sub_740_47_n_133 & sub_740_47_n_30) | ~(sub_740_47_n_133 | sub_740_47_n_30));
 assign sub_740_47_n_138 = ~(sub_740_47_n_135 & ~sub_740_47_n_41);
 assign T_14_32_ = ~sub_740_47_n_136;
 assign sub_740_47_n_136 = ~(sub_740_47_n_125 & ~sub_740_47_n_102);
 assign sub_740_47_n_135 = ~(sub_740_47_n_34 & ~sub_740_47_n_92);
 assign sub_740_47_n_134 = ~(sub_740_47_n_127 & ~sub_740_47_n_4);
 assign sub_740_47_n_133 = ~(sub_740_47_n_126 & ~sub_740_47_n_1);
 assign T_14_16_ = ((sub_740_47_n_124 & sub_740_47_n_83) | ~(sub_740_47_n_124 | sub_740_47_n_83));
 assign T_14_12_ = ((sub_740_47_n_123 & sub_740_47_n_27) | ~(sub_740_47_n_123 | sub_740_47_n_27));
 assign T_14_10_ = ((sub_740_47_n_35 & sub_740_47_n_28) | ~(sub_740_47_n_35 | sub_740_47_n_28));
 assign T_14_9_ = ((sub_740_47_n_122 & sub_740_47_n_23) | ~(sub_740_47_n_122 | sub_740_47_n_23));
 assign T_14_7_ = ((sub_740_47_n_20 & sub_740_47_n_19) | ~(sub_740_47_n_20 | sub_740_47_n_19));
 assign sub_740_47_n_127 = ~(sub_740_47_n_123 & ~sub_740_47_n_64);
 assign sub_740_47_n_126 = ~(sub_740_47_n_35 & ~sub_740_47_n_61);
 assign sub_740_47_n_125 = ~(sub_740_47_n_124 & ~sub_740_47_n_37);
 assign sub_740_47_n_124 = ~(sub_740_47_n_115 & sub_740_47_n_36);
 assign sub_740_47_n_123 = ~(sub_740_47_n_118 & ~sub_740_47_n_101);
 assign sub_740_47_n_122 = ~(sub_740_47_n_117 & ~sub_740_47_n_3);
 assign T_14_6_ = ((sub_740_47_n_113 & sub_740_47_n_16) | ~(sub_740_47_n_113 | sub_740_47_n_16));
 assign T_14_5_ = ~((sub_740_47_n_15 | sub_740_47_n_13) & ~(sub_740_47_n_15 & sub_740_47_n_13));
 assign T_14_8_ = ((sub_740_47_n_114 & sub_740_47_n_17) | ~(sub_740_47_n_114 | sub_740_47_n_17));
 assign sub_740_47_n_118 = ~(sub_740_47_n_114 & ~sub_740_47_n_95);
 assign sub_740_47_n_117 = ~(sub_740_47_n_114 & ~sub_740_47_n_52);
 assign sub_740_47_n_116 = ~(sub_740_47_n_113 & ~sub_740_47_n_51);
 assign sub_740_47_n_115 = ~(sub_740_47_n_114 & sub_740_47_n_99);
 assign sub_740_47_n_114 = ~(sub_740_47_n_109 & sub_740_47_n_100);
 assign sub_740_47_n_113 = ~(sub_740_47_n_31 & ~sub_740_47_n_90);
 assign T_14_4_ = ~((sub_740_47_n_108 | sub_740_47_n_25) & ~(sub_740_47_n_108 & sub_740_47_n_25));
 assign T_14_3_ = ((sub_740_47_n_24 & sub_740_47_n_26) | ~(sub_740_47_n_24 | sub_740_47_n_26));
 assign sub_740_47_n_110 = ~(sub_740_47_n_108 & ~sub_740_47_n_62);
 assign sub_740_47_n_109 = ~(sub_740_47_n_108 & ~sub_740_47_n_94);
 assign sub_740_47_n_108 = ~(sub_740_47_n_105 & sub_740_47_n_87);
 assign T_14_2_ = ~((sub_740_47_n_104 | sub_740_47_n_29) & ~(sub_740_47_n_104 & sub_740_47_n_29));
 assign sub_740_47_n_106 = ~(sub_740_47_n_104 & ~sub_740_47_n_65);
 assign sub_740_47_n_105 = ~(sub_740_47_n_104 & sub_740_47_n_81);
 assign sub_740_47_n_104 = ((n_1189 & R_15_0_) | ((R_15_0_ & sub_740_47_n_46) | (sub_740_47_n_46 & n_1189)));
 assign T_14_1_ = (R_15_0_ ^ (sub_740_47_n_46 ^ n_1189));
 assign sub_740_47_n_102 = ~(sub_740_47_n_98 | (sub_740_47_n_69 & (sub_740_47_n_56 | sub_740_47_n_66)));
 assign sub_740_47_n_101 = ~(sub_740_47_n_93 & (sub_740_47_n_96 | sub_740_47_n_79));
 assign sub_740_47_n_100 = ~(sub_740_47_n_89 | (sub_740_47_n_90 & sub_740_47_n_84));
 assign sub_740_47_n_99 = ~(sub_740_47_n_95 | sub_740_47_n_97);
 assign sub_740_47_n_98 = ~(sub_740_47_n_72 & (sub_740_47_n_71 & (sub_740_47_n_74 & sub_740_47_n_75)));
 assign sub_740_47_n_94 = ~(sub_740_47_n_76 & sub_740_47_n_84);
 assign sub_740_47_n_93 = ~(sub_740_47_n_68 | (sub_740_47_n_1 & sub_740_47_n_59));
 assign sub_740_47_n_97 = ~(sub_740_47_n_86 & sub_740_47_n_77);
 assign sub_740_47_n_96 = ~(sub_740_47_n_10 | (sub_740_47_n_3 & sub_740_47_n_55));
 assign sub_740_47_n_95 = ~(sub_740_47_n_82 & sub_740_47_n_78);
 assign sub_740_47_n_92 = ~sub_740_47_n_91;
 assign sub_740_47_n_89 = ~(sub_740_47_n_8 & (sub_740_47_n_42 | sub_740_47_n_53));
 assign sub_740_47_n_88 = ~(sub_740_47_n_11 | (sub_740_47_n_40 & sub_740_47_n_50));
 assign sub_740_47_n_87 = ~(sub_740_47_n_80 | ~sub_740_47_n_6);
 assign sub_740_47_n_91 = ~(sub_740_47_n_70 | (~sub_740_47_n_39 & sub_740_47_n_4));
 assign sub_740_47_n_90 = ~(sub_740_47_n_2 & (sub_740_47_n_5 | sub_740_47_n_38));
 assign sub_740_47_n_81 = ~(sub_740_47_n_65 | sub_740_47_n_63);
 assign sub_740_47_n_80 = ~(sub_740_47_n_43 | sub_740_47_n_63);
 assign sub_740_47_n_86 = ~(sub_740_47_n_64 | sub_740_47_n_39);
 assign sub_740_47_n_85 = ~(sub_740_47_n_69 & sub_740_47_n_67);
 assign sub_740_47_n_84 = ~(sub_740_47_n_51 | sub_740_47_n_53);
 assign sub_740_47_n_83 = ~(sub_740_47_n_56 & sub_740_47_n_0);
 assign sub_740_47_n_79 = ~(sub_740_47_n_60 & sub_740_47_n_59);
 assign sub_740_47_n_78 = ~(sub_740_47_n_61 | sub_740_47_n_58);
 assign sub_740_47_n_82 = ~(sub_740_47_n_52 | sub_740_47_n_54);
 assign sub_740_47_n_75 = ~(n_1361 | (n_830 | n_1273));
 assign sub_740_47_n_74 = ~(n_1086 | (n_1242 | n_1297));
 assign T_14_0_ = ~(sub_740_47_n_57 & (~{in2[14]} | {in1[0]}));
 assign sub_740_47_n_72 = ~(n_1031 | (n_1302 | (n_1212 | n_1366)));
 assign sub_740_47_n_71 = ~(n_1177 | (n_1292 | (n_1059 | n_1371)));
 assign sub_740_47_n_77 = ~(sub_740_47_n_41 | sub_740_47_n_49);
 assign sub_740_47_n_76 = ~(sub_740_47_n_62 | sub_740_47_n_38);
 assign sub_740_47_n_70 = ~sub_740_47_n_7;
 assign sub_740_47_n_67 = ~sub_740_47_n_66;
 assign sub_740_47_n_60 = ~sub_740_47_n_61;
 assign sub_740_47_n_58 = ~sub_740_47_n_59;
 assign sub_740_47_n_69 = ~(R_15_16_ & ~n_1172);
 assign sub_740_47_n_68 = ~(n_1065 | sub_740_47_n_47);
 assign sub_740_47_n_66 = ~(R_15_16_ | ~n_1172);
 assign sub_740_47_n_65 = ~(R_15_1_ | ~n_1101);
 assign sub_740_47_n_64 = ~(R_15_11_ | ~n_1026);
 assign sub_740_47_n_63 = ~(R_15_2_ | ~n_1113);
 assign sub_740_47_n_62 = ~(R_15_3_ | ~n_1340);
 assign sub_740_47_n_43 = ~(R_15_1_ & ~n_1101);
 assign sub_740_47_n_61 = ~(R_15_9_ | ~n_1345);
 assign sub_740_47_n_59 = ~(sub_740_47_n_47 & ~sub_740_47_n_48);
 assign sub_740_47_n_57 = ~({in1[0]} & ~{in2[14]});
 assign sub_740_47_n_55 = ~sub_740_47_n_54;
 assign sub_740_47_n_50 = ~sub_740_47_n_49;
 assign sub_740_47_n_40 = ~sub_740_47_n_9;
 assign sub_740_47_n_56 = ~(sub_740_47_n_45 & R_15_15_);
 assign sub_740_47_n_54 = ~(R_15_8_ | ~n_1162);
 assign sub_740_47_n_42 = ~(R_15_5_ & ~n_1096);
 assign sub_740_47_n_53 = ~(R_15_6_ | ~n_1167);
 assign sub_740_47_n_41 = ~(R_15_13_ | ~n_1182);
 assign sub_740_47_n_52 = ~(R_15_7_ | ~n_1217);
 assign sub_740_47_n_51 = ~(R_15_5_ | ~n_1096);
 assign sub_740_47_n_49 = ~(R_15_14_ | ~n_1091);
 assign sub_740_47_n_48 = ~n_1065;
 assign sub_740_47_n_47 = ~R_15_10_;
 assign sub_740_47_n_46 = ~n_1350;
 assign sub_740_47_n_45 = ~n_1136;
 assign sub_740_47_n_39 = ~(R_15_12_ | ~n_1259);
 assign sub_740_47_n_38 = ~(R_15_4_ | ~n_1049);
 assign sub_740_47_n_37 = ~(sub_740_47_n_67 & (sub_740_47_n_0 & ~sub_740_47_n_98));
 assign sub_740_47_n_36 = ~(sub_740_47_n_32 | (~sub_740_47_n_97 & sub_740_47_n_101));
 assign sub_740_47_n_35 = ~(sub_740_47_n_33 & sub_740_47_n_96);
 assign sub_740_47_n_34 = ~(sub_740_47_n_123 & sub_740_47_n_86);
 assign sub_740_47_n_33 = ~(sub_740_47_n_114 & sub_740_47_n_82);
 assign sub_740_47_n_32 = ~(sub_740_47_n_88 & (~sub_740_47_n_77 | sub_740_47_n_91));
 assign sub_740_47_n_31 = ~(sub_740_47_n_108 & sub_740_47_n_76);
 assign sub_740_47_n_30 = ~(sub_740_47_n_59 & ~sub_740_47_n_68);
 assign sub_740_47_n_29 = ~(sub_740_47_n_43 & ~sub_740_47_n_65);
 assign sub_740_47_n_28 = ~(sub_740_47_n_60 & ~sub_740_47_n_1);
 assign sub_740_47_n_27 = (sub_740_47_n_4 | sub_740_47_n_64);
 assign sub_740_47_n_26 = ~(sub_740_47_n_6 & ~sub_740_47_n_63);
 assign sub_740_47_n_25 = ~(sub_740_47_n_5 & ~sub_740_47_n_62);
 assign sub_740_47_n_24 = ~(sub_740_47_n_106 & sub_740_47_n_43);
 assign sub_740_47_n_23 = ~(sub_740_47_n_55 & ~sub_740_47_n_10);
 assign sub_740_47_n_22 = ~(sub_740_47_n_50 & ~sub_740_47_n_11);
 assign sub_740_47_n_21 = ~(sub_740_47_n_14 & sub_740_47_n_56);
 assign sub_740_47_n_20 = ~(sub_740_47_n_116 & sub_740_47_n_42);
 assign sub_740_47_n_19 = ~(sub_740_47_n_8 & ~sub_740_47_n_53);
 assign sub_740_47_n_18 = ~(sub_740_47_n_9 & ~sub_740_47_n_41);
 assign sub_740_47_n_17 = (sub_740_47_n_3 | sub_740_47_n_52);
 assign sub_740_47_n_16 = ~(sub_740_47_n_42 & ~sub_740_47_n_51);
 assign sub_740_47_n_15 = ~(sub_740_47_n_110 & sub_740_47_n_5);
 assign sub_740_47_n_14 = ~(sub_740_47_n_124 & sub_740_47_n_0);
 assign sub_740_47_n_13 = ~(sub_740_47_n_2 & ~sub_740_47_n_38);
 assign sub_740_47_n_12 = ~(sub_740_47_n_7 & ~sub_740_47_n_39);
 assign sub_740_47_n_11 = ~(n_1091 | ~R_15_14_);
 assign sub_740_47_n_10 = ~(n_1162 | ~R_15_8_);
 assign sub_740_47_n_9 = ~(R_15_13_ & ~n_1182);
 assign sub_740_47_n_8 = ~(R_15_6_ & ~n_1167);
 assign sub_740_47_n_7 = ~(R_15_12_ & ~n_1259);
 assign sub_740_47_n_6 = ~(R_15_2_ & ~n_1113);
 assign sub_740_47_n_5 = ~(R_15_3_ & ~n_1340);
 assign sub_740_47_n_4 = ~(n_1026 | ~R_15_11_);
 assign sub_740_47_n_3 = ~(n_1217 | ~R_15_7_);
 assign sub_740_47_n_2 = ~(R_15_4_ & ~n_1049);
 assign sub_740_47_n_1 = ~(n_1345 | ~R_15_9_);
 assign sub_740_47_n_0 = (R_15_15_ | sub_740_47_n_45);
 assign T_13_15_ = ~((sub_770_46_n_31 | sub_770_46_n_21) & ~(sub_770_46_n_31 & sub_770_46_n_21));
 assign T_13_18_ = ((sub_770_46_n_145 & sub_770_46_n_20) | ~(sub_770_46_n_145 | sub_770_46_n_20));
 assign T_13_17_ = ((sub_770_46_n_144 & sub_770_46_n_90) | ~(sub_770_46_n_144 | sub_770_46_n_90));
 assign T_13_14_ = ((sub_770_46_n_34 & sub_770_46_n_86) | ~(sub_770_46_n_34 | sub_770_46_n_86));
 assign T_13_13_ = ((sub_770_46_n_143 & sub_770_46_n_23) | ~(sub_770_46_n_143 | sub_770_46_n_23));
 assign T_13_11_ = ((sub_770_46_n_141 & sub_770_46_n_74) | ~(sub_770_46_n_141 | sub_770_46_n_74));
 assign T_13_32_ = ~sub_770_46_n_142;
 assign sub_770_46_n_142 = ~(sub_770_46_n_136 & ~sub_770_46_n_112);
 assign sub_770_46_n_145 = ~(sub_770_46_n_103 & (~sub_770_46_n_85 | sub_770_46_n_134));
 assign sub_770_46_n_144 = ~(sub_770_46_n_62 & (~sub_770_46_n_48 | sub_770_46_n_134));
 assign sub_770_46_n_143 = ~(sub_770_46_n_64 & (~sub_770_46_n_0 | sub_770_46_n_28));
 assign T_13_10_ = ~((sub_770_46_n_132 | sub_770_46_n_81) & ~(sub_770_46_n_132 & sub_770_46_n_81));
 assign T_13_12_ = ~((sub_770_46_n_135 | sub_770_46_n_75) & ~(sub_770_46_n_135 & sub_770_46_n_75));
 assign T_13_16_ = ((sub_770_46_n_40 & sub_770_46_n_88) | ~(sub_770_46_n_40 | sub_770_46_n_88));
 assign T_13_7_ = ((sub_770_46_n_129 & sub_770_46_n_79) | ~(sub_770_46_n_129 | sub_770_46_n_79));
 assign sub_770_46_n_141 = ~(sub_770_46_n_37 & (~sub_770_46_n_2 | sub_770_46_n_131));
 assign sub_770_46_n_136 = ~(sub_770_46_n_133 & ~sub_770_46_n_29);
 assign sub_770_46_n_135 = ~sub_770_46_n_28;
 assign sub_770_46_n_40 = ~sub_770_46_n_134;
 assign sub_770_46_n_134 = ~sub_770_46_n_133;
 assign sub_770_46_n_133 = ~(sub_770_46_n_115 & (sub_770_46_n_125 | sub_770_46_n_109));
 assign sub_770_46_n_132 = ~sub_770_46_n_131;
 assign sub_770_46_n_131 = ~(sub_770_46_n_100 | (~sub_770_46_n_80 & sub_770_46_n_126));
 assign sub_770_46_n_130 = ~(sub_770_46_n_50 & (~sub_770_46_n_5 | sub_770_46_n_127));
 assign sub_770_46_n_129 = ~(sub_770_46_n_35 & (~sub_770_46_n_12 | sub_770_46_n_124));
 assign T_13_8_ = ((sub_770_46_n_127 & sub_770_46_n_18) | ~(sub_770_46_n_127 | sub_770_46_n_18));
 assign sub_770_46_n_127 = ~sub_770_46_n_126;
 assign sub_770_46_n_126 = ~sub_770_46_n_125;
 assign sub_770_46_n_125 = ~(sub_770_46_n_110 | (sub_770_46_n_104 & sub_770_46_n_118));
 assign sub_770_46_n_124 = ~(sub_770_46_n_102 | (~sub_770_46_n_95 & sub_770_46_n_118));
 assign sub_770_46_n_123 = ~(sub_770_46_n_60 & (~sub_770_46_n_7 | sub_770_46_n_119));
 assign T_13_4_ = ((sub_770_46_n_119 & sub_770_46_n_24) | ~(sub_770_46_n_119 | sub_770_46_n_24));
 assign T_13_3_ = ((sub_770_46_n_120 & sub_770_46_n_77) | ~(sub_770_46_n_120 | sub_770_46_n_77));
 assign sub_770_46_n_120 = ~(sub_770_46_n_6 | (~sub_770_46_n_63 & sub_770_46_n_114));
 assign sub_770_46_n_119 = ~sub_770_46_n_118;
 assign sub_770_46_n_118 = ~(sub_770_46_n_116 & sub_770_46_n_17);
 assign T_13_2_ = ~((sub_770_46_n_114 | sub_770_46_n_22) & ~(sub_770_46_n_114 & sub_770_46_n_22));
 assign sub_770_46_n_116 = ~(sub_770_46_n_114 & sub_770_46_n_83);
 assign sub_770_46_n_115 = ~(sub_770_46_n_33 | (sub_770_46_n_111 & sub_770_46_n_26));
 assign sub_770_46_n_114 = ((n_1153 & n_979) | ((n_979 & n_1354) | (n_1354 & n_1153)));
 assign T_13_1_ = (n_979 ^ (n_1354 ^ n_1153));
 assign sub_770_46_n_112 = ~(sub_770_46_n_108 | (sub_770_46_n_82 & (sub_770_46_n_103 | sub_770_46_n_94)));
 assign sub_770_46_n_111 = ~(sub_770_46_n_98 & (sub_770_46_n_99 | sub_770_46_n_87));
 assign sub_770_46_n_110 = ~(sub_770_46_n_97 & (sub_770_46_n_101 | sub_770_46_n_78));
 assign sub_770_46_n_109 = ~(sub_770_46_n_107 & sub_770_46_n_26);
 assign sub_770_46_n_108 = ~(sub_770_46_n_73 & (sub_770_46_n_72 & (sub_770_46_n_69 & sub_770_46_n_70)));
 assign sub_770_46_n_106 = ~sub_770_46_n_105;
 assign sub_770_46_n_104 = ~(sub_770_46_n_95 | sub_770_46_n_78);
 assign sub_770_46_n_107 = ~(sub_770_46_n_80 | sub_770_46_n_87);
 assign sub_770_46_n_105 = ~(sub_770_46_n_68 & (sub_770_46_n_64 | sub_770_46_n_65));
 assign sub_770_46_n_102 = ~sub_770_46_n_101;
 assign sub_770_46_n_100 = ~sub_770_46_n_99;
 assign sub_770_46_n_98 = ~(sub_770_46_n_67 | (sub_770_46_n_57 & sub_770_46_n_15));
 assign sub_770_46_n_97 = ~(sub_770_46_n_54 | (sub_770_46_n_51 & sub_770_46_n_8));
 assign sub_770_46_n_96 = ~(sub_770_46_n_1 & (sub_770_46_n_9 | sub_770_46_n_61));
 assign sub_770_46_n_103 = ~(sub_770_46_n_84 | ~sub_770_46_n_53);
 assign sub_770_46_n_101 = ~(sub_770_46_n_66 | (sub_770_46_n_4 & sub_770_46_n_16));
 assign sub_770_46_n_99 = ~(sub_770_46_n_11 | (sub_770_46_n_49 & sub_770_46_n_10));
 assign sub_770_46_n_94 = ~sub_770_46_n_3;
 assign sub_770_46_n_93 = ~sub_770_46_n_92;
 assign sub_770_46_n_84 = ~(sub_770_46_n_62 | ~sub_770_46_n_13);
 assign sub_770_46_n_83 = ~(sub_770_46_n_63 | sub_770_46_n_52);
 assign sub_770_46_n_82 = ~(sub_770_46_n_14 & ~n_1303);
 assign sub_770_46_n_95 = ~(sub_770_46_n_7 & sub_770_46_n_16);
 assign sub_770_46_n_92 = ~(sub_770_46_n_0 & ~sub_770_46_n_65);
 assign sub_770_46_n_91 = ~(sub_770_46_n_35 & sub_770_46_n_12);
 assign sub_770_46_n_90 = ~(sub_770_46_n_53 & sub_770_46_n_13);
 assign sub_770_46_n_89 = ~(sub_770_46_n_38 & sub_770_46_n_16);
 assign sub_770_46_n_88 = ~(sub_770_46_n_62 & sub_770_46_n_48);
 assign sub_770_46_n_87 = ~(sub_770_46_n_2 & sub_770_46_n_15);
 assign sub_770_46_n_86 = ~(sub_770_46_n_9 & sub_770_46_n_59);
 assign sub_770_46_n_85 = ~(sub_770_46_n_47 | ~sub_770_46_n_13);
 assign sub_770_46_n_73 = ~(n_1213 | (n_1367 | n_1178));
 assign sub_770_46_n_72 = ~(n_1293 | (n_1060 | n_1372));
 assign T_13_0_ = ~(sub_770_46_n_56 & (~{in2[13]} | {in1[0]}));
 assign sub_770_46_n_70 = ~(n_1362 | (n_831 | n_1274));
 assign sub_770_46_n_69 = ~(n_1087 | (n_1243 | n_1298));
 assign sub_770_46_n_81 = ~(sub_770_46_n_37 & sub_770_46_n_2);
 assign sub_770_46_n_80 = ~(sub_770_46_n_5 & sub_770_46_n_10);
 assign sub_770_46_n_79 = ~(sub_770_46_n_36 & sub_770_46_n_8);
 assign sub_770_46_n_78 = ~(sub_770_46_n_12 & sub_770_46_n_8);
 assign sub_770_46_n_77 = ~(sub_770_46_n_32 | sub_770_46_n_52);
 assign sub_770_46_n_76 = ~(sub_770_46_n_58 | sub_770_46_n_61);
 assign sub_770_46_n_75 = ~(sub_770_46_n_64 & sub_770_46_n_0);
 assign sub_770_46_n_74 = ~(sub_770_46_n_39 & sub_770_46_n_15);
 assign sub_770_46_n_67 = ~sub_770_46_n_39;
 assign sub_770_46_n_66 = ~sub_770_46_n_38;
 assign sub_770_46_n_60 = ~sub_770_46_n_4;
 assign sub_770_46_n_59 = ~sub_770_46_n_58;
 assign sub_770_46_n_57 = ~sub_770_46_n_37;
 assign sub_770_46_n_68 = ~(n_973 & ~n_1260);
 assign sub_770_46_n_39 = ~(sub_770_46_n_45 & n_984);
 assign sub_770_46_n_38 = ~(n_985 & ~n_1050);
 assign sub_770_46_n_65 = ~(n_973 | ~n_1260);
 assign sub_770_46_n_64 = ~(sub_770_46_n_43 & R_14_11_);
 assign sub_770_46_n_63 = ~(n_966 | ~n_1102);
 assign sub_770_46_n_62 = ~(R_14_15_ & ~n_1137);
 assign sub_770_46_n_61 = ~(n_986 | ~n_1092);
 assign sub_770_46_n_58 = ~(n_972 | ~n_1183);
 assign sub_770_46_n_37 = ~(n_970 & ~n_1346);
 assign sub_770_46_n_56 = ~({in1[0]} & ~{in2[13]});
 assign sub_770_46_n_54 = ~sub_770_46_n_36;
 assign sub_770_46_n_51 = ~sub_770_46_n_35;
 assign sub_770_46_n_50 = ~sub_770_46_n_49;
 assign sub_770_46_n_48 = ~sub_770_46_n_47;
 assign sub_770_46_n_55 = ~(R_14_17_ | ~n_1032);
 assign sub_770_46_n_36 = ~(sub_770_46_n_46 & n_977);
 assign sub_770_46_n_53 = ~(n_980 & ~n_1173);
 assign sub_770_46_n_52 = ~(n_969 | ~n_1114);
 assign sub_770_46_n_35 = ~(n_971 & ~n_1097);
 assign sub_770_46_n_49 = ~(n_1218 | sub_770_46_n_44);
 assign sub_770_46_n_47 = ~(R_14_15_ | ~n_1137);
 assign sub_770_46_n_46 = ~n_1168;
 assign sub_770_46_n_45 = ~n_1066;
 assign sub_770_46_n_44 = ~n_978;
 assign sub_770_46_n_43 = ~n_1027;
 assign sub_770_46_n_42 = ~n_1350;
 assign sub_770_46_n_34 = ~(sub_770_46_n_106 & (~sub_770_46_n_93 | sub_770_46_n_28));
 assign sub_770_46_n_33 = (sub_770_46_n_96 | (sub_770_46_n_105 & sub_770_46_n_76));
 assign sub_770_46_n_32 = ~(n_1114 | ~n_969);
 assign sub_770_46_n_31 = ~(sub_770_46_n_9 & ~(sub_770_46_n_59 & sub_770_46_n_34));
 assign T_13_6_ = (sub_770_46_n_124 ^ sub_770_46_n_91);
 assign sub_770_46_n_29 = ~(sub_770_46_n_3 & (sub_770_46_n_85 & ~sub_770_46_n_108));
 assign sub_770_46_n_28 = ~(sub_770_46_n_111 | (sub_770_46_n_107 & sub_770_46_n_126));
 assign T_13_5_ = ~(sub_770_46_n_123 ^ sub_770_46_n_89);
 assign sub_770_46_n_26 = ~(sub_770_46_n_92 | ~sub_770_46_n_76);
 assign T_13_9_ = ~(sub_770_46_n_130 ^ sub_770_46_n_19);
 assign sub_770_46_n_24 = ~(sub_770_46_n_4 | ~sub_770_46_n_7);
 assign sub_770_46_n_23 = ~(sub_770_46_n_68 & ~sub_770_46_n_65);
 assign sub_770_46_n_22 = (sub_770_46_n_6 | sub_770_46_n_63);
 assign sub_770_46_n_21 = ~(sub_770_46_n_1 & ~sub_770_46_n_61);
 assign sub_770_46_n_20 = (sub_770_46_n_14 | sub_770_46_n_55);
 assign sub_770_46_n_19 = ~(sub_770_46_n_10 & ~sub_770_46_n_11);
 assign sub_770_46_n_18 = ~(sub_770_46_n_49 | ~sub_770_46_n_5);
 assign sub_770_46_n_17 = ~(sub_770_46_n_32 | (~sub_770_46_n_52 & sub_770_46_n_6));
 assign sub_770_46_n_16 = ~(n_1050 & ~n_985);
 assign sub_770_46_n_15 = (n_984 | sub_770_46_n_45);
 assign sub_770_46_n_14 = ~(n_1032 | ~R_14_17_);
 assign sub_770_46_n_13 = ~(n_1173 & ~n_980);
 assign sub_770_46_n_12 = ~(n_1097 & ~n_971);
 assign sub_770_46_n_11 = ~(n_1163 | ~n_968);
 assign sub_770_46_n_10 = ~(n_1163 & ~n_968);
 assign sub_770_46_n_9 = ~(n_972 & ~n_1183);
 assign sub_770_46_n_8 = (n_977 | sub_770_46_n_46);
 assign sub_770_46_n_7 = ~(n_1341 & ~n_967);
 assign sub_770_46_n_6 = ~(n_1102 | ~n_966);
 assign sub_770_46_n_5 = ~(sub_770_46_n_44 & n_1218);
 assign sub_770_46_n_4 = ~(n_1341 | ~n_967);
 assign sub_770_46_n_3 = ~(sub_770_46_n_55 | n_1303);
 assign sub_770_46_n_2 = ~(n_1346 & ~n_970);
 assign sub_770_46_n_1 = ~(n_986 & ~n_1092);
 assign sub_770_46_n_0 = (R_14_11_ | sub_770_46_n_43);
 assign T_12_15_ = ~(sub_800_45_n_167 & sub_800_45_n_169);
 assign T_12_19_ = ((sub_800_45_n_168 & sub_800_45_n_20) | ~(sub_800_45_n_168 | sub_800_45_n_20));
 assign sub_800_45_n_169 = ~(sub_800_45_n_16 & (sub_800_45_n_161 | sub_800_45_n_57));
 assign sub_800_45_n_168 = ~(sub_800_45_n_66 | (sub_800_45_n_155 & sub_800_45_n_63));
 assign sub_800_45_n_167 = ~(sub_800_45_n_160 & (~sub_800_45_n_16 & ~sub_800_45_n_57));
 assign T_12_18_ = ((sub_800_45_n_155 & sub_800_45_n_88) | ~(sub_800_45_n_155 | sub_800_45_n_88));
 assign T_12_17_ = ((sub_800_45_n_158 & sub_800_45_n_24) | ~(sub_800_45_n_158 | sub_800_45_n_24));
 assign T_12_14_ = ~((sub_800_45_n_156 | sub_800_45_n_91) & ~(sub_800_45_n_156 & sub_800_45_n_91));
 assign T_12_13_ = ((sub_800_45_n_159 & sub_800_45_n_25) | ~(sub_800_45_n_159 | sub_800_45_n_25));
 assign T_12_11_ = ((sub_800_45_n_153 & sub_800_45_n_26) | ~(sub_800_45_n_153 | sub_800_45_n_26));
 assign sub_800_45_n_161 = ~(sub_800_45_n_157 | ~sub_800_45_n_64);
 assign sub_800_45_n_160 = ~(sub_800_45_n_156 & ~sub_800_45_n_29);
 assign sub_800_45_n_157 = ~sub_800_45_n_156;
 assign T_12_32_ = ~(sub_800_45_n_146 | ~sub_800_45_n_118);
 assign sub_800_45_n_159 = ~(sub_800_45_n_68 | (~sub_800_45_n_65 & sub_800_45_n_145));
 assign sub_800_45_n_158 = ~(sub_800_45_n_52 | (~sub_800_45_n_45 & sub_800_45_n_143));
 assign sub_800_45_n_156 = ~(sub_800_45_n_147 & ~sub_800_45_n_104);
 assign sub_800_45_n_155 = ~(sub_800_45_n_107 & (sub_800_45_n_142 | sub_800_45_n_77));
 assign T_12_10_ = ((sub_800_45_n_141 & sub_800_45_n_83) | ~(sub_800_45_n_141 | sub_800_45_n_83));
 assign T_12_12_ = ~((sub_800_45_n_145 | sub_800_45_n_22) & ~(sub_800_45_n_145 & sub_800_45_n_22));
 assign T_12_16_ = ((sub_800_45_n_144 & sub_800_45_n_85) | ~(sub_800_45_n_144 | sub_800_45_n_85));
 assign T_12_9_ = ((sub_800_45_n_139 & sub_800_45_n_18) | ~(sub_800_45_n_139 | sub_800_45_n_18));
 assign T_12_7_ = ~((sub_800_45_n_138 | sub_800_45_n_81) & ~(sub_800_45_n_138 & sub_800_45_n_81));
 assign sub_800_45_n_153 = ~(sub_800_45_n_44 | (~sub_800_45_n_41 & sub_800_45_n_140));
 assign sub_800_45_n_147 = ~(sub_800_45_n_145 & ~sub_800_45_n_90);
 assign sub_800_45_n_146 = ~(sub_800_45_n_142 | ~sub_800_45_n_117);
 assign sub_800_45_n_145 = ~(sub_800_45_n_134 & ~sub_800_45_n_115);
 assign sub_800_45_n_144 = ~sub_800_45_n_143;
 assign sub_800_45_n_143 = ~sub_800_45_n_142;
 assign sub_800_45_n_142 = ~(sub_800_45_n_132 | sub_800_45_n_120);
 assign sub_800_45_n_141 = ~sub_800_45_n_140;
 assign sub_800_45_n_140 = ~(sub_800_45_n_133 & ~sub_800_45_n_98);
 assign sub_800_45_n_139 = ~(sub_800_45_n_42 | (~sub_800_45_n_54 & sub_800_45_n_131));
 assign sub_800_45_n_138 = ~(sub_800_45_n_30 & (~sub_800_45_n_14 | sub_800_45_n_129));
 assign T_12_6_ = ((sub_800_45_n_129 & sub_800_45_n_15) | ~(sub_800_45_n_129 | sub_800_45_n_15));
 assign T_12_5_ = ~((sub_800_45_n_128 | sub_800_45_n_19) & ~(sub_800_45_n_128 & sub_800_45_n_19));
 assign T_12_8_ = ~((sub_800_45_n_131 | sub_800_45_n_17) & ~(sub_800_45_n_131 & sub_800_45_n_17));
 assign sub_800_45_n_134 = ~(sub_800_45_n_131 & ~sub_800_45_n_105);
 assign sub_800_45_n_133 = ~(sub_800_45_n_131 & ~sub_800_45_n_79);
 assign sub_800_45_n_132 = ~(sub_800_45_n_130 | ~sub_800_45_n_109);
 assign sub_800_45_n_131 = ~sub_800_45_n_130;
 assign sub_800_45_n_130 = ~(sub_800_45_n_113 | (sub_800_45_n_123 & sub_800_45_n_102));
 assign sub_800_45_n_129 = ~(sub_800_45_n_100 | (~sub_800_45_n_93 & sub_800_45_n_123));
 assign sub_800_45_n_128 = ~(sub_800_45_n_47 & (~sub_800_45_n_13 | sub_800_45_n_124));
 assign T_12_4_ = ((sub_800_45_n_124 & sub_800_45_n_21) | ~(sub_800_45_n_124 | sub_800_45_n_21));
 assign T_12_3_ = ((sub_800_45_n_125 & sub_800_45_n_86) | ~(sub_800_45_n_125 | sub_800_45_n_86));
 assign sub_800_45_n_125 = ~(sub_800_45_n_121 & ~sub_800_45_n_69);
 assign sub_800_45_n_124 = ~sub_800_45_n_123;
 assign sub_800_45_n_123 = ~(sub_800_45_n_101 & (sub_800_45_n_111 | sub_800_45_n_82));
 assign T_12_2_ = ~((sub_800_45_n_119 | sub_800_45_n_23) & ~(sub_800_45_n_119 & sub_800_45_n_23));
 assign sub_800_45_n_121 = ~(sub_800_45_n_119 & ~sub_800_45_n_49);
 assign sub_800_45_n_120 = ~(sub_800_45_n_112 & (sub_800_45_n_114 | sub_800_45_n_103));
 assign sub_800_45_n_119 = ~sub_800_45_n_111;
 assign sub_800_45_n_118 = ~(sub_800_45_n_108 & (sub_800_45_n_95 | (sub_800_45_n_106 & sub_800_45_n_92)));
 assign sub_800_45_n_117 = ~(sub_800_45_n_116 | sub_800_45_n_77);
 assign sub_800_45_n_116 = ~(sub_800_45_n_108 & sub_800_45_n_92);
 assign sub_800_45_n_115 = ~sub_800_45_n_114;
 assign sub_800_45_n_114 = ~(sub_800_45_n_97 | (sub_800_45_n_98 & sub_800_45_n_84));
 assign sub_800_45_n_113 = ~(sub_800_45_n_94 & (sub_800_45_n_99 | sub_800_45_n_80));
 assign sub_800_45_n_112 = ~(sub_800_45_n_96 | (sub_800_45_n_104 & sub_800_45_n_87));
 assign sub_800_45_n_111 = ~((n_1268 & R_13_0_) | ((R_13_0_ & sub_800_45_n_35) | (sub_800_45_n_35 & n_1268)));
 assign T_12_1_ = ~(R_13_0_ ^ (n_1351 ^ n_1268));
 assign sub_800_45_n_109 = ~(sub_800_45_n_105 | sub_800_45_n_103);
 assign sub_800_45_n_108 = (sub_800_45_n_75 & (sub_800_45_n_73 & (sub_800_45_n_76 & sub_800_45_n_74)));
 assign sub_800_45_n_107 = ~sub_800_45_n_106;
 assign sub_800_45_n_102 = ~(sub_800_45_n_93 | sub_800_45_n_80);
 assign sub_800_45_n_101 = ~(sub_800_45_n_71 | (sub_800_45_n_69 & sub_800_45_n_8));
 assign sub_800_45_n_106 = ~(sub_800_45_n_70 & (~sub_800_45_n_60 | sub_800_45_n_51));
 assign sub_800_45_n_105 = ~(sub_800_45_n_78 & sub_800_45_n_84);
 assign sub_800_45_n_104 = ~(sub_800_45_n_4 & (sub_800_45_n_67 | sub_800_45_n_59));
 assign sub_800_45_n_103 = ~(sub_800_45_n_89 & sub_800_45_n_87);
 assign sub_800_45_n_100 = ~sub_800_45_n_99;
 assign sub_800_45_n_97 = ~(sub_800_45_n_12 & (sub_800_45_n_43 | sub_800_45_n_27));
 assign sub_800_45_n_96 = ~(sub_800_45_n_3 & (sub_800_45_n_56 | sub_800_45_n_50));
 assign sub_800_45_n_95 = ~(sub_800_45_n_1 & (sub_800_45_n_2 | sub_800_45_n_53));
 assign sub_800_45_n_94 = ~(sub_800_45_n_55 | (sub_800_45_n_31 & sub_800_45_n_7));
 assign sub_800_45_n_99 = ~(sub_800_45_n_10 | (sub_800_45_n_46 & sub_800_45_n_11));
 assign sub_800_45_n_98 = ~(sub_800_45_n_5 & (sub_800_45_n_0 | sub_800_45_n_48));
 assign sub_800_45_n_90 = ~sub_800_45_n_89;
 assign sub_800_45_n_82 = ~(sub_800_45_n_9 & sub_800_45_n_8);
 assign sub_800_45_n_93 = ~(sub_800_45_n_13 & sub_800_45_n_11);
 assign sub_800_45_n_92 = ~(sub_800_45_n_62 | sub_800_45_n_53);
 assign sub_800_45_n_91 = ~(sub_800_45_n_56 & sub_800_45_n_64);
 assign sub_800_45_n_89 = ~(sub_800_45_n_65 | sub_800_45_n_59);
 assign sub_800_45_n_88 = ~(sub_800_45_n_2 & sub_800_45_n_63);
 assign sub_800_45_n_87 = ~(sub_800_45_n_29 | sub_800_45_n_50);
 assign sub_800_45_n_86 = ~(sub_800_45_n_32 & sub_800_45_n_8);
 assign sub_800_45_n_85 = ~(sub_800_45_n_52 | sub_800_45_n_45);
 assign sub_800_45_n_84 = ~(sub_800_45_n_40 | sub_800_45_n_27);
 assign sub_800_45_n_83 = ~(sub_800_45_n_44 | sub_800_45_n_41);
 assign sub_800_45_n_79 = ~sub_800_45_n_78;
 assign sub_800_45_n_76 = ~(n_1087 | (n_1243 | n_1298));
 assign sub_800_45_n_75 = ~(n_1213 | (n_1367 | n_1178));
 assign sub_800_45_n_74 = ~(n_1362 | (n_831 | n_1274));
 assign sub_800_45_n_73 = ~(n_1293 | (n_1060 | n_1372));
 assign T_12_0_ = ~(sub_800_45_n_58 & (~{in2[12]} | {in1[0]}));
 assign sub_800_45_n_81 = ~(sub_800_45_n_28 & sub_800_45_n_7);
 assign sub_800_45_n_80 = ~(sub_800_45_n_14 & sub_800_45_n_7);
 assign sub_800_45_n_78 = ~(sub_800_45_n_54 | sub_800_45_n_48);
 assign sub_800_45_n_77 = ~(sub_800_45_n_6 & ~sub_800_45_n_61);
 assign sub_800_45_n_71 = ~sub_800_45_n_32;
 assign sub_800_45_n_31 = ~sub_800_45_n_30;
 assign sub_800_45_n_68 = ~sub_800_45_n_67;
 assign sub_800_45_n_66 = ~sub_800_45_n_2;
 assign sub_800_45_n_64 = ~sub_800_45_n_29;
 assign sub_800_45_n_63 = ~sub_800_45_n_62;
 assign sub_800_45_n_61 = ~sub_800_45_n_60;
 assign sub_800_45_n_57 = ~sub_800_45_n_56;
 assign sub_800_45_n_32 = ~(R_13_2_ & ~n_1114);
 assign sub_800_45_n_70 = ~(sub_800_45_n_38 & R_13_16_);
 assign sub_800_45_n_30 = ~(R_13_5_ & ~n_1097);
 assign sub_800_45_n_69 = ~(n_1102 | sub_800_45_n_39);
 assign sub_800_45_n_67 = ~(R_13_11_ & ~n_1027);
 assign sub_800_45_n_65 = ~(R_13_11_ | ~n_1027);
 assign sub_800_45_n_29 = ~(R_13_13_ | ~n_1183);
 assign sub_800_45_n_62 = ~(R_13_17_ | ~n_1032);
 assign sub_800_45_n_60 = ~(sub_800_45_n_34 & ~sub_800_45_n_38);
 assign sub_800_45_n_59 = ~(R_13_12_ | ~n_1260);
 assign sub_800_45_n_58 = ~({in1[0]} & ~{in2[12]});
 assign sub_800_45_n_56 = ~(R_13_13_ & ~n_1183);
 assign sub_800_45_n_55 = ~sub_800_45_n_28;
 assign sub_800_45_n_52 = ~sub_800_45_n_51;
 assign sub_800_45_n_49 = ~sub_800_45_n_9;
 assign sub_800_45_n_47 = ~sub_800_45_n_46;
 assign sub_800_45_n_45 = ~sub_800_45_n_6;
 assign sub_800_45_n_44 = ~sub_800_45_n_43;
 assign sub_800_45_n_42 = ~sub_800_45_n_0;
 assign sub_800_45_n_28 = ~(sub_800_45_n_36 & R_13_6_);
 assign sub_800_45_n_54 = ~(R_13_7_ | ~n_1218);
 assign sub_800_45_n_53 = ~(R_13_18_ | ~n_1303);
 assign sub_800_45_n_51 = ~(R_13_15_ & ~n_1137);
 assign sub_800_45_n_50 = ~(R_13_14_ | ~n_1092);
 assign sub_800_45_n_48 = ~(R_13_8_ | ~n_1163);
 assign sub_800_45_n_46 = ~(n_1341 | sub_800_45_n_37);
 assign sub_800_45_n_43 = ~(R_13_9_ & ~n_1346);
 assign sub_800_45_n_40 = ~(R_13_9_ | ~n_1346);
 assign sub_800_45_n_41 = ~(R_13_9_ | ~n_1346);
 assign sub_800_45_n_39 = ~R_13_1_;
 assign sub_800_45_n_38 = ~n_1173;
 assign sub_800_45_n_37 = ~R_13_3_;
 assign sub_800_45_n_36 = ~n_1168;
 assign sub_800_45_n_35 = ~n_1351;
 assign sub_800_45_n_34 = ~R_13_16_;
 assign sub_800_45_n_27 = ~(R_13_10_ | ~n_1066);
 assign sub_800_45_n_26 = ~(sub_800_45_n_27 | ~sub_800_45_n_12);
 assign sub_800_45_n_25 = ~(sub_800_45_n_59 | ~sub_800_45_n_4);
 assign sub_800_45_n_24 = ~(sub_800_45_n_61 | ~sub_800_45_n_70);
 assign sub_800_45_n_23 = (sub_800_45_n_69 | sub_800_45_n_49);
 assign sub_800_45_n_22 = ~(sub_800_45_n_67 & ~sub_800_45_n_65);
 assign sub_800_45_n_21 = (sub_800_45_n_47 & sub_800_45_n_13);
 assign sub_800_45_n_20 = ~(sub_800_45_n_53 | ~sub_800_45_n_1);
 assign sub_800_45_n_19 = ~(sub_800_45_n_11 & ~sub_800_45_n_10);
 assign sub_800_45_n_18 = ~(sub_800_45_n_48 | ~sub_800_45_n_5);
 assign sub_800_45_n_17 = ~(sub_800_45_n_0 & ~sub_800_45_n_54);
 assign sub_800_45_n_16 = ~(sub_800_45_n_3 & ~sub_800_45_n_50);
 assign sub_800_45_n_15 = ~(sub_800_45_n_31 | ~sub_800_45_n_14);
 assign sub_800_45_n_14 = ~(n_1097 & ~R_13_5_);
 assign sub_800_45_n_13 = ~(sub_800_45_n_37 & n_1341);
 assign sub_800_45_n_12 = ~(R_13_10_ & ~n_1066);
 assign sub_800_45_n_11 = ~(n_1050 & ~R_13_4_);
 assign sub_800_45_n_10 = ~(n_1050 | ~R_13_4_);
 assign sub_800_45_n_9 = ~(sub_800_45_n_39 & n_1102);
 assign sub_800_45_n_8 = ~(n_1114 & ~R_13_2_);
 assign sub_800_45_n_7 = (R_13_6_ | sub_800_45_n_36);
 assign sub_800_45_n_6 = ~(n_1137 & ~R_13_15_);
 assign sub_800_45_n_5 = ~(R_13_8_ & ~n_1163);
 assign sub_800_45_n_4 = ~(R_13_12_ & ~n_1260);
 assign sub_800_45_n_3 = ~(R_13_14_ & ~n_1092);
 assign sub_800_45_n_2 = ~(R_13_17_ & ~n_1032);
 assign sub_800_45_n_1 = ~(R_13_18_ & ~n_1303);
 assign sub_800_45_n_0 = ~(R_13_7_ & ~n_1218);
 assign T_11_19_ = ((sub_830_44_n_182 & sub_830_44_n_26) | ~(sub_830_44_n_182 | sub_830_44_n_26));
 assign T_11_15_ = ((sub_830_44_n_23 & sub_830_44_n_27) | ~(sub_830_44_n_23 | sub_830_44_n_27));
 assign sub_830_44_n_182 = ~(sub_830_44_n_16 | ~sub_830_44_n_6);
 assign T_11_20_ = ((sub_830_44_n_34 & sub_830_44_n_28) | ~(sub_830_44_n_34 | sub_830_44_n_28));
 assign T_11_18_ = ((sub_830_44_n_172 & sub_830_44_n_107) | ~(sub_830_44_n_172 | sub_830_44_n_107));
 assign T_11_17_ = ((sub_830_44_n_174 & sub_830_44_n_22) | ~(sub_830_44_n_174 | sub_830_44_n_22));
 assign T_11_14_ = ((sub_830_44_n_173 & sub_830_44_n_93) | ~(sub_830_44_n_173 | sub_830_44_n_93));
 assign T_11_13_ = ((sub_830_44_n_18 & sub_830_44_n_102) | ~(sub_830_44_n_18 | sub_830_44_n_102));
 assign T_11_11_ = ((sub_830_44_n_15 & sub_830_44_n_19) | ~(sub_830_44_n_15 | sub_830_44_n_19));
 assign T_11_32_ = ~sub_830_44_n_171;
 assign sub_830_44_n_171 = ~(sub_830_44_n_161 & sub_830_44_n_147);
 assign sub_830_44_n_174 = ~(sub_830_44_n_163 | ~sub_830_44_n_39);
 assign sub_830_44_n_173 = ~(sub_830_44_n_162 & ~sub_830_44_n_119);
 assign sub_830_44_n_172 = ~(sub_830_44_n_164 | ~sub_830_44_n_120);
 assign T_11_9_ = ~((sub_830_44_n_157 | sub_830_44_n_21) & ~(sub_830_44_n_157 & sub_830_44_n_21));
 assign T_11_10_ = ~((sub_830_44_n_33 | sub_830_44_n_24) & ~(sub_830_44_n_33 & sub_830_44_n_24));
 assign T_11_12_ = ((sub_830_44_n_160 & sub_830_44_n_101) | ~(sub_830_44_n_160 | sub_830_44_n_101));
 assign T_11_7_ = ((sub_830_44_n_17 & sub_830_44_n_97) | ~(sub_830_44_n_17 | sub_830_44_n_97));
 assign T_11_16_ = ((sub_830_44_n_159 & sub_830_44_n_20) | ~(sub_830_44_n_159 | sub_830_44_n_20));
 assign sub_830_44_n_165 = ~(sub_830_44_n_159 | ~sub_830_44_n_126);
 assign sub_830_44_n_164 = ~(sub_830_44_n_159 | ~sub_830_44_n_95);
 assign sub_830_44_n_163 = ~(sub_830_44_n_159 | ~sub_830_44_n_9);
 assign sub_830_44_n_162 = ~(sub_830_44_n_160 & ~sub_830_44_n_108);
 assign sub_830_44_n_161 = ~(sub_830_44_n_158 & ~sub_830_44_n_138);
 assign sub_830_44_n_160 = ~(sub_830_44_n_137 & (~sub_830_44_n_125 | sub_830_44_n_153));
 assign sub_830_44_n_159 = ~sub_830_44_n_158;
 assign sub_830_44_n_158 = ~(sub_830_44_n_141 & (sub_830_44_n_46 | sub_830_44_n_131));
 assign sub_830_44_n_157 = ~(sub_830_44_n_69 & (~sub_830_44_n_8 | sub_830_44_n_46));
 assign T_11_6_ = ((sub_830_44_n_152 & sub_830_44_n_109) | ~(sub_830_44_n_152 | sub_830_44_n_109));
 assign T_11_8_ = ((sub_830_44_n_47 & sub_830_44_n_106) | ~(sub_830_44_n_47 | sub_830_44_n_106));
 assign sub_830_44_n_154 = ~(sub_830_44_n_47 & ~sub_830_44_n_99);
 assign sub_830_44_n_153 = ~sub_830_44_n_47;
 assign sub_830_44_n_47 = ~sub_830_44_n_46;
 assign sub_830_44_n_46 = ~(sub_830_44_n_133 | (sub_830_44_n_144 & sub_830_44_n_122));
 assign sub_830_44_n_152 = ~sub_830_44_n_151;
 assign sub_830_44_n_151 = ~(sub_830_44_n_124 | (~sub_830_44_n_113 & sub_830_44_n_144));
 assign sub_830_44_n_150 = ~(sub_830_44_n_78 & (sub_830_44_n_145 | sub_830_44_n_85));
 assign T_11_4_ = ~((sub_830_44_n_145 | sub_830_44_n_105) & ~(sub_830_44_n_145 & sub_830_44_n_105));
 assign T_11_3_ = ((sub_830_44_n_146 & sub_830_44_n_30) | ~(sub_830_44_n_146 | sub_830_44_n_30));
 assign sub_830_44_n_147 = ~(sub_830_44_n_127 & (sub_830_44_n_31 | (sub_830_44_n_134 & sub_830_44_n_130)));
 assign sub_830_44_n_146 = ~(sub_830_44_n_77 | (sub_830_44_n_140 & sub_830_44_n_83));
 assign sub_830_44_n_145 = ~sub_830_44_n_144;
 assign sub_830_44_n_144 = ~(sub_830_44_n_142 & sub_830_44_n_117);
 assign T_11_2_ = ~((sub_830_44_n_140 | sub_830_44_n_111) & ~(sub_830_44_n_140 & sub_830_44_n_111));
 assign sub_830_44_n_142 = ~(sub_830_44_n_140 & sub_830_44_n_103);
 assign sub_830_44_n_141 = ~(sub_830_44_n_135 | (sub_830_44_n_136 & sub_830_44_n_128));
 assign sub_830_44_n_140 = ((n_1074 & R_12_0_) | ((R_12_0_ & sub_830_44_n_49) | (sub_830_44_n_49 & n_1074)));
 assign T_11_1_ = (R_12_0_ ^ (sub_830_44_n_49 ^ n_1074));
 assign sub_830_44_n_138 = ~(sub_830_44_n_132 & sub_830_44_n_126);
 assign sub_830_44_n_137 = ~sub_830_44_n_136;
 assign sub_830_44_n_136 = ~(sub_830_44_n_118 & (sub_830_44_n_121 | sub_830_44_n_100));
 assign sub_830_44_n_135 = ~(sub_830_44_n_116 & (sub_830_44_n_25 | sub_830_44_n_112));
 assign sub_830_44_n_134 = ~(sub_830_44_n_114 & (~sub_830_44_n_110 | sub_830_44_n_120));
 assign sub_830_44_n_133 = ~(sub_830_44_n_115 & (sub_830_44_n_123 | sub_830_44_n_98));
 assign sub_830_44_n_132 = ~(sub_830_44_n_129 | ~sub_830_44_n_127);
 assign sub_830_44_n_131 = ~(sub_830_44_n_125 & sub_830_44_n_128);
 assign sub_830_44_n_130 = ~sub_830_44_n_129;
 assign sub_830_44_n_124 = ~sub_830_44_n_123;
 assign sub_830_44_n_122 = ~(sub_830_44_n_113 | sub_830_44_n_98);
 assign sub_830_44_n_129 = ~(sub_830_44_n_96 & sub_830_44_n_10);
 assign sub_830_44_n_128 = ~(sub_830_44_n_108 | sub_830_44_n_112);
 assign sub_830_44_n_127 = (sub_830_44_n_89 & sub_830_44_n_92);
 assign sub_830_44_n_126 = ~(sub_830_44_n_94 | ~sub_830_44_n_110);
 assign sub_830_44_n_125 = ~(sub_830_44_n_99 | sub_830_44_n_100);
 assign sub_830_44_n_123 = ~(sub_830_44_n_12 | (sub_830_44_n_7 & sub_830_44_n_11));
 assign sub_830_44_n_119 = ~sub_830_44_n_25;
 assign sub_830_44_n_118 = ~(sub_830_44_n_87 | (sub_830_44_n_74 & sub_830_44_n_2));
 assign sub_830_44_n_117 = ~(sub_830_44_n_104 | ~sub_830_44_n_88);
 assign sub_830_44_n_116 = ~(sub_830_44_n_35 | (sub_830_44_n_45 & sub_830_44_n_84));
 assign sub_830_44_n_115 = ~(sub_830_44_n_71 | (sub_830_44_n_64 & sub_830_44_n_81));
 assign sub_830_44_n_114 = ~(sub_830_44_n_36 | (sub_830_44_n_76 & sub_830_44_n_80));
 assign sub_830_44_n_121 = ~(sub_830_44_n_70 | (sub_830_44_n_68 & sub_830_44_n_13));
 assign sub_830_44_n_120 = ~(sub_830_44_n_90 | ~sub_830_44_n_4);
 assign sub_830_44_n_104 = ~(sub_830_44_n_43 | sub_830_44_n_65);
 assign sub_830_44_n_103 = ~(sub_830_44_n_82 | sub_830_44_n_65);
 assign sub_830_44_n_113 = ~(sub_830_44_n_14 & sub_830_44_n_11);
 assign sub_830_44_n_112 = ~(sub_830_44_n_73 & sub_830_44_n_84);
 assign sub_830_44_n_111 = ~(sub_830_44_n_43 & sub_830_44_n_83);
 assign sub_830_44_n_110 = ~(sub_830_44_n_38 | sub_830_44_n_79);
 assign sub_830_44_n_109 = ~(sub_830_44_n_37 & sub_830_44_n_66);
 assign sub_830_44_n_108 = ~(sub_830_44_n_5 & ~sub_830_44_n_75);
 assign sub_830_44_n_107 = ~(sub_830_44_n_76 | sub_830_44_n_38);
 assign sub_830_44_n_106 = ~(sub_830_44_n_69 & sub_830_44_n_8);
 assign sub_830_44_n_105 = ~(sub_830_44_n_7 | sub_830_44_n_85);
 assign sub_830_44_n_95 = ~sub_830_44_n_94;
 assign sub_830_44_n_92 = ~(n_1298 | (n_1362 | (n_831 | n_1274)));
 assign T_11_0_ = ~(sub_830_44_n_72 & (~{in2[11]} | {in1[0]}));
 assign sub_830_44_n_90 = ~(sub_830_44_n_39 | ~sub_830_44_n_3);
 assign sub_830_44_n_89 = ~(n_1060 | (n_1372 | (n_1087 | n_1243)));
 assign sub_830_44_n_102 = ~(sub_830_44_n_0 | sub_830_44_n_75);
 assign sub_830_44_n_101 = ~(sub_830_44_n_41 & sub_830_44_n_5);
 assign sub_830_44_n_100 = ~(sub_830_44_n_1 & sub_830_44_n_2);
 assign sub_830_44_n_99 = ~(sub_830_44_n_8 & sub_830_44_n_13);
 assign sub_830_44_n_98 = ~(sub_830_44_n_66 & sub_830_44_n_81);
 assign sub_830_44_n_97 = ~(sub_830_44_n_40 & sub_830_44_n_81);
 assign sub_830_44_n_96 = ~(n_1178 | (n_1293 | n_1367));
 assign sub_830_44_n_94 = ~(sub_830_44_n_9 & ~sub_830_44_n_67);
 assign sub_830_44_n_93 = ~(sub_830_44_n_44 & sub_830_44_n_73);
 assign sub_830_44_n_45 = ~sub_830_44_n_44;
 assign sub_830_44_n_85 = ~sub_830_44_n_14;
 assign sub_830_44_n_83 = ~sub_830_44_n_82;
 assign sub_830_44_n_80 = ~sub_830_44_n_79;
 assign sub_830_44_n_78 = ~sub_830_44_n_7;
 assign sub_830_44_n_77 = ~sub_830_44_n_43;
 assign sub_830_44_n_76 = ~sub_830_44_n_6;
 assign sub_830_44_n_42 = ~sub_830_44_n_41;
 assign sub_830_44_n_88 = ~(sub_830_44_n_52 & R_12_2_);
 assign sub_830_44_n_87 = ~(n_1066 | sub_830_44_n_62);
 assign sub_830_44_n_86 = ~(R_12_19_ & ~n_1213);
 assign sub_830_44_n_44 = ~(R_12_13_ & ~n_1183);
 assign sub_830_44_n_84 = ~(sub_830_44_n_54 & ~sub_830_44_n_58);
 assign sub_830_44_n_82 = ~(R_12_1_ | ~n_1102);
 assign sub_830_44_n_81 = ~(sub_830_44_n_57 & ~sub_830_44_n_53);
 assign sub_830_44_n_79 = ~(R_12_18_ | ~n_1303);
 assign sub_830_44_n_43 = ~(R_12_1_ & ~n_1102);
 assign sub_830_44_n_75 = ~(R_12_12_ | ~n_1260);
 assign sub_830_44_n_41 = ~(R_12_11_ & ~n_1027);
 assign sub_830_44_n_74 = ~(n_1346 | sub_830_44_n_60);
 assign sub_830_44_n_73 = ~(sub_830_44_n_63 & ~sub_830_44_n_50);
 assign sub_830_44_n_72 = ~({in1[0]} & ~{in2[11]});
 assign sub_830_44_n_71 = ~sub_830_44_n_40;
 assign sub_830_44_n_69 = ~sub_830_44_n_68;
 assign sub_830_44_n_67 = ~sub_830_44_n_3;
 assign sub_830_44_n_64 = ~sub_830_44_n_37;
 assign sub_830_44_n_40 = ~(sub_830_44_n_53 & R_12_6_);
 assign sub_830_44_n_70 = ~(n_1163 | sub_830_44_n_51);
 assign sub_830_44_n_39 = ~(R_12_15_ & ~n_1137);
 assign sub_830_44_n_68 = ~(n_1218 | sub_830_44_n_56);
 assign sub_830_44_n_66 = ~(sub_830_44_n_61 & ~sub_830_44_n_59);
 assign sub_830_44_n_65 = ~(R_12_2_ | ~n_1114);
 assign sub_830_44_n_38 = ~(R_12_17_ | ~n_1032);
 assign sub_830_44_n_37 = ~(sub_830_44_n_59 & R_12_5_);
 assign sub_830_44_n_63 = ~R_12_13_;
 assign sub_830_44_n_62 = ~R_12_10_;
 assign sub_830_44_n_61 = ~R_12_5_;
 assign sub_830_44_n_60 = ~R_12_9_;
 assign sub_830_44_n_59 = ~n_1097;
 assign sub_830_44_n_58 = ~n_1092;
 assign sub_830_44_n_57 = ~R_12_6_;
 assign sub_830_44_n_56 = ~R_12_7_;
 assign sub_830_44_n_55 = ~R_12_16_;
 assign sub_830_44_n_54 = ~R_12_14_;
 assign sub_830_44_n_53 = ~n_1168;
 assign sub_830_44_n_52 = ~n_1114;
 assign sub_830_44_n_51 = ~R_12_8_;
 assign sub_830_44_n_50 = ~n_1183;
 assign sub_830_44_n_49 = ~n_1351;
 assign sub_830_44_n_36 = ~(n_1303 | ~R_12_18_);
 assign sub_830_44_n_35 = (sub_830_44_n_58 & R_12_14_);
 assign sub_830_44_n_34 = ~(sub_830_44_n_165 | sub_830_44_n_134);
 assign sub_830_44_n_33 = ~(sub_830_44_n_154 & sub_830_44_n_121);
 assign T_11_5_ = ~(sub_830_44_n_150 ^ sub_830_44_n_29);
 assign sub_830_44_n_31 = ~(sub_830_44_n_86 | ~sub_830_44_n_96);
 assign sub_830_44_n_30 = ~(sub_830_44_n_65 | ~sub_830_44_n_88);
 assign sub_830_44_n_29 = ~(sub_830_44_n_11 & ~sub_830_44_n_12);
 assign sub_830_44_n_28 = (sub_830_44_n_86 & sub_830_44_n_10);
 assign sub_830_44_n_27 = ~(sub_830_44_n_35 | ~sub_830_44_n_84);
 assign sub_830_44_n_26 = ~(sub_830_44_n_36 | ~sub_830_44_n_80);
 assign sub_830_44_n_25 = ~(sub_830_44_n_0 | (~sub_830_44_n_75 & sub_830_44_n_42));
 assign sub_830_44_n_24 = ~(sub_830_44_n_1 & ~sub_830_44_n_74);
 assign sub_830_44_n_23 = ~(sub_830_44_n_45 | (sub_830_44_n_73 & sub_830_44_n_173));
 assign sub_830_44_n_22 = ~(sub_830_44_n_67 | ~sub_830_44_n_4);
 assign sub_830_44_n_21 = ~(sub_830_44_n_13 & ~sub_830_44_n_70);
 assign sub_830_44_n_20 = (sub_830_44_n_39 & sub_830_44_n_9);
 assign sub_830_44_n_19 = ~(sub_830_44_n_87 | ~sub_830_44_n_2);
 assign sub_830_44_n_18 = ~(sub_830_44_n_42 | (sub_830_44_n_5 & sub_830_44_n_160));
 assign sub_830_44_n_17 = ~(sub_830_44_n_37 & (~sub_830_44_n_66 | sub_830_44_n_151));
 assign sub_830_44_n_16 = ~(sub_830_44_n_172 | sub_830_44_n_38);
 assign sub_830_44_n_15 = ~(sub_830_44_n_74 | (sub_830_44_n_1 & sub_830_44_n_33));
 assign sub_830_44_n_14 = ~(n_1341 & ~R_12_3_);
 assign sub_830_44_n_13 = ~(sub_830_44_n_51 & n_1163);
 assign sub_830_44_n_12 = ~(n_1050 | ~R_12_4_);
 assign sub_830_44_n_11 = ~(n_1050 & ~R_12_4_);
 assign sub_830_44_n_10 = ~(n_1213 & ~R_12_19_);
 assign sub_830_44_n_9 = ~(n_1137 & ~R_12_15_);
 assign sub_830_44_n_8 = ~(sub_830_44_n_56 & n_1218);
 assign sub_830_44_n_7 = ~(n_1341 | ~R_12_3_);
 assign sub_830_44_n_6 = ~(R_12_17_ & ~n_1032);
 assign sub_830_44_n_5 = ~(n_1027 & ~R_12_11_);
 assign sub_830_44_n_4 = (sub_830_44_n_55 | n_1173);
 assign sub_830_44_n_3 = ~(sub_830_44_n_55 & n_1173);
 assign sub_830_44_n_2 = ~(sub_830_44_n_62 & n_1066);
 assign sub_830_44_n_1 = ~(sub_830_44_n_60 & n_1346);
 assign sub_830_44_n_0 = ~(n_1260 | ~R_12_12_);
 assign T_10_21_ = ((sub_860_43_n_20 & sub_860_43_n_18) | ~(sub_860_43_n_20 | sub_860_43_n_18));
 assign T_10_19_ = ((sub_860_43_n_23 & sub_860_43_n_101) | ~(sub_860_43_n_23 | sub_860_43_n_101));
 assign T_10_15_ = ((sub_860_43_n_176 & sub_860_43_n_21) | ~(sub_860_43_n_176 | sub_860_43_n_21));
 assign sub_860_43_n_176 = ~(sub_860_43_n_80 | (~sub_860_43_n_73 & sub_860_43_n_166));
 assign T_10_20_ = ((sub_860_43_n_165 & sub_860_43_n_19) | ~(sub_860_43_n_165 | sub_860_43_n_19));
 assign T_10_18_ = ((sub_860_43_n_167 & sub_860_43_n_99) | ~(sub_860_43_n_167 | sub_860_43_n_99));
 assign T_10_17_ = ((sub_860_43_n_169 & sub_860_43_n_25) | ~(sub_860_43_n_169 | sub_860_43_n_25));
 assign T_10_14_ = ((sub_860_43_n_166 & sub_860_43_n_24) | ~(sub_860_43_n_166 | sub_860_43_n_24));
 assign T_10_13_ = ((sub_860_43_n_168 & sub_860_43_n_22) | ~(sub_860_43_n_168 | sub_860_43_n_22));
 assign T_10_11_ = ((sub_860_43_n_163 & sub_860_43_n_30) | ~(sub_860_43_n_163 | sub_860_43_n_30));
 assign T_10_32_ = ~(sub_860_43_n_141 | sub_860_43_n_158);
 assign sub_860_43_n_169 = ~(sub_860_43_n_76 | (~sub_860_43_n_57 & sub_860_43_n_157));
 assign sub_860_43_n_168 = ~(sub_860_43_n_52 | (sub_860_43_n_35 & sub_860_43_n_65));
 assign sub_860_43_n_167 = ~(sub_860_43_n_115 | (~sub_860_43_n_104 & sub_860_43_n_157));
 assign sub_860_43_n_166 = ~(sub_860_43_n_32 & ~sub_860_43_n_112);
 assign sub_860_43_n_165 = ~(sub_860_43_n_131 | (~sub_860_43_n_121 & sub_860_43_n_157));
 assign T_10_9_ = ((sub_860_43_n_155 & sub_860_43_n_15) | ~(sub_860_43_n_155 | sub_860_43_n_15));
 assign T_10_10_ = ((sub_860_43_n_43 & sub_860_43_n_90) | ~(sub_860_43_n_43 | sub_860_43_n_90));
 assign T_10_12_ = ~((sub_860_43_n_35 | sub_860_43_n_95) & ~(sub_860_43_n_35 & sub_860_43_n_95));
 assign T_10_7_ = ((sub_860_43_n_154 & sub_860_43_n_92) | ~(sub_860_43_n_154 | sub_860_43_n_92));
 assign sub_860_43_n_163 = ~(sub_860_43_n_56 | (~sub_860_43_n_61 & sub_860_43_n_156));
 assign sub_860_43_n_158 = ~(sub_860_43_n_44 | ~sub_860_43_n_133);
 assign sub_860_43_n_157 = ~sub_860_43_n_44;
 assign sub_860_43_n_44 = ~(sub_860_43_n_149 | sub_860_43_n_137);
 assign sub_860_43_n_43 = ~sub_860_43_n_156;
 assign sub_860_43_n_156 = ~(sub_860_43_n_31 & ~sub_860_43_n_113);
 assign sub_860_43_n_155 = ~(sub_860_43_n_8 & (~sub_860_43_n_54 | sub_860_43_n_146));
 assign sub_860_43_n_154 = ~(sub_860_43_n_40 & (~sub_860_43_n_7 | sub_860_43_n_147));
 assign T_10_6_ = ~((sub_860_43_n_147 | sub_860_43_n_16) & ~(sub_860_43_n_147 & sub_860_43_n_16));
 assign T_10_5_ = ~((sub_860_43_n_148 | sub_860_43_n_28) & ~(sub_860_43_n_148 & sub_860_43_n_28));
 assign T_10_8_ = ~((sub_860_43_n_145 | sub_860_43_n_93) & ~(sub_860_43_n_145 & sub_860_43_n_93));
 assign sub_860_43_n_150 = ~(sub_860_43_n_145 & ~sub_860_43_n_120);
 assign sub_860_43_n_149 = ~(sub_860_43_n_146 | ~sub_860_43_n_125);
 assign sub_860_43_n_148 = ~(sub_860_43_n_142 | ~sub_860_43_n_60);
 assign sub_860_43_n_147 = ~(sub_860_43_n_33 | ~sub_860_43_n_122);
 assign sub_860_43_n_145 = ~sub_860_43_n_146;
 assign sub_860_43_n_146 = ~(sub_860_43_n_128 | (sub_860_43_n_116 & sub_860_43_n_139));
 assign T_10_4_ = ((sub_860_43_n_140 & sub_860_43_n_29) | ~(sub_860_43_n_140 | sub_860_43_n_29));
 assign T_10_3_ = ((sub_860_43_n_26 & sub_860_43_n_17) | ~(sub_860_43_n_26 | sub_860_43_n_17));
 assign sub_860_43_n_142 = ~(sub_860_43_n_140 | ~sub_860_43_n_5);
 assign sub_860_43_n_141 = ~(sub_860_43_n_117 | (~sub_860_43_n_124 & sub_860_43_n_135));
 assign sub_860_43_n_140 = ~sub_860_43_n_139;
 assign sub_860_43_n_139 = ~(sub_860_43_n_136 & sub_860_43_n_107);
 assign T_10_2_ = ~((sub_860_43_n_134 | sub_860_43_n_27) & ~(sub_860_43_n_134 & sub_860_43_n_27));
 assign sub_860_43_n_137 = ~(sub_860_43_n_130 & (sub_860_43_n_129 | sub_860_43_n_123));
 assign sub_860_43_n_136 = ~(sub_860_43_n_14 & (sub_860_43_n_13 & sub_860_43_n_134));
 assign sub_860_43_n_135 = ~(sub_860_43_n_131 & ~sub_860_43_n_119);
 assign sub_860_43_n_134 = ~(sub_860_43_n_126 & (sub_860_43_n_127 & sub_860_43_n_67));
 assign sub_860_43_n_133 = ~(sub_860_43_n_34 | sub_860_43_n_121);
 assign T_10_1_ = ~((sub_860_43_n_91 | n_1210) & ~(sub_860_43_n_91 & n_1210));
 assign sub_860_43_n_131 = ~(sub_860_43_n_110 & (~sub_860_43_n_100 | sub_860_43_n_114));
 assign sub_860_43_n_130 = ~(sub_860_43_n_111 | (sub_860_43_n_112 & sub_860_43_n_105));
 assign sub_860_43_n_129 = ~(sub_860_43_n_108 | (sub_860_43_n_113 & sub_860_43_n_97));
 assign sub_860_43_n_128 = ~(sub_860_43_n_109 & (sub_860_43_n_122 | sub_860_43_n_96));
 assign sub_860_43_n_127 = ~(n_1210 & R_11_0_);
 assign sub_860_43_n_126 = ~(n_1210 & ~n_1351);
 assign sub_860_43_n_125 = ~(sub_860_43_n_120 | sub_860_43_n_123);
 assign sub_860_43_n_124 = ~(sub_860_43_n_69 | (sub_860_43_n_1 & (sub_860_43_n_39 | sub_860_43_n_63)));
 assign sub_860_43_n_119 = ~sub_860_43_n_118;
 assign sub_860_43_n_116 = ~(sub_860_43_n_106 | sub_860_43_n_96);
 assign sub_860_43_n_123 = ~(sub_860_43_n_102 & sub_860_43_n_105);
 assign sub_860_43_n_122 = ~(sub_860_43_n_37 | (sub_860_43_n_59 & sub_860_43_n_11));
 assign sub_860_43_n_121 = ~(sub_860_43_n_103 & sub_860_43_n_100);
 assign sub_860_43_n_120 = ~(sub_860_43_n_94 & sub_860_43_n_97);
 assign sub_860_43_n_118 = ~(sub_860_43_n_69 | (sub_860_43_n_63 | sub_860_43_n_66));
 assign sub_860_43_n_117 = ~(sub_860_43_n_87 & sub_860_43_n_88);
 assign sub_860_43_n_115 = ~sub_860_43_n_114;
 assign sub_860_43_n_111 = ~(sub_860_43_n_6 & (sub_860_43_n_2 | sub_860_43_n_82));
 assign sub_860_43_n_110 = ~(sub_860_43_n_84 | (sub_860_43_n_81 & sub_860_43_n_78));
 assign sub_860_43_n_109 = ~(sub_860_43_n_85 | (sub_860_43_n_79 & sub_860_43_n_9));
 assign sub_860_43_n_108 = ~(sub_860_43_n_4 & (sub_860_43_n_55 | sub_860_43_n_71));
 assign sub_860_43_n_107 = ~(sub_860_43_n_38 | (sub_860_43_n_83 & sub_860_43_n_13));
 assign sub_860_43_n_114 = ~(sub_860_43_n_89 | ~sub_860_43_n_68);
 assign sub_860_43_n_113 = ~(sub_860_43_n_12 & (sub_860_43_n_8 | sub_860_43_n_58));
 assign sub_860_43_n_112 = ~(sub_860_43_n_3 & (sub_860_43_n_51 | sub_860_43_n_62));
 assign sub_860_43_n_104 = ~sub_860_43_n_103;
 assign sub_860_43_n_106 = ~(sub_860_43_n_5 & sub_860_43_n_11);
 assign sub_860_43_n_105 = ~(sub_860_43_n_73 | sub_860_43_n_82);
 assign sub_860_43_n_103 = ~(sub_860_43_n_57 | ~sub_860_43_n_74);
 assign sub_860_43_n_102 = ~(sub_860_43_n_64 | sub_860_43_n_62);
 assign sub_860_43_n_101 = ~(sub_860_43_n_10 & sub_860_43_n_78);
 assign sub_860_43_n_100 = ~(sub_860_43_n_72 | sub_860_43_n_77);
 assign sub_860_43_n_99 = ~(sub_860_43_n_81 | sub_860_43_n_72);
 assign sub_860_43_n_98 = ~(sub_860_43_n_76 | sub_860_43_n_57);
 assign sub_860_43_n_97 = ~(sub_860_43_n_61 | sub_860_43_n_71);
 assign sub_860_43_n_89 = ~(sub_860_43_n_75 | ~sub_860_43_n_74);
 assign sub_860_43_n_88 = ~(n_1298 | (n_1362 | (n_831 | n_1274)));
 assign sub_860_43_n_87 = ~(n_1060 | (n_1372 | (n_1087 | n_1243)));
 assign T_10_0_ = ~(sub_860_43_n_70 & (~{in2[10]} | {in1[0]}));
 assign sub_860_43_n_96 = ~(sub_860_43_n_7 & sub_860_43_n_9);
 assign sub_860_43_n_95 = ~(sub_860_43_n_51 & sub_860_43_n_65);
 assign sub_860_43_n_94 = ~(sub_860_43_n_53 | sub_860_43_n_58);
 assign sub_860_43_n_93 = ~(sub_860_43_n_8 & sub_860_43_n_54);
 assign sub_860_43_n_92 = ~(sub_860_43_n_42 & sub_860_43_n_9);
 assign sub_860_43_n_91 = ~(sub_860_43_n_67 & sub_860_43_n_0);
 assign sub_860_43_n_90 = ~(sub_860_43_n_56 | sub_860_43_n_61);
 assign sub_860_43_n_85 = ~sub_860_43_n_42;
 assign sub_860_43_n_84 = ~sub_860_43_n_10;
 assign sub_860_43_n_81 = ~sub_860_43_n_41;
 assign sub_860_43_n_80 = ~sub_860_43_n_2;
 assign sub_860_43_n_79 = ~sub_860_43_n_40;
 assign sub_860_43_n_78 = ~sub_860_43_n_77;
 assign sub_860_43_n_76 = ~sub_860_43_n_75;
 assign sub_860_43_n_42 = ~(sub_860_43_n_49 & R_11_6_);
 assign sub_860_43_n_83 = ~(n_1102 | sub_860_43_n_47);
 assign sub_860_43_n_82 = ~(R_11_14_ | ~n_1092);
 assign sub_860_43_n_41 = ~(R_11_17_ & ~n_1032);
 assign sub_860_43_n_40 = ~(R_11_5_ & ~n_1097);
 assign sub_860_43_n_77 = ~(R_11_18_ | ~n_1303);
 assign sub_860_43_n_75 = ~(R_11_15_ & ~n_1137);
 assign sub_860_43_n_74 = ~(sub_860_43_n_46 & ~sub_860_43_n_50);
 assign sub_860_43_n_73 = ~(R_11_13_ | ~n_1183);
 assign sub_860_43_n_72 = ~(R_11_17_ | ~n_1032);
 assign sub_860_43_n_71 = ~(R_11_10_ | ~n_1066);
 assign sub_860_43_n_70 = ~({in1[0]} & ~{in2[10]});
 assign sub_860_43_n_65 = ~sub_860_43_n_64;
 assign sub_860_43_n_60 = ~sub_860_43_n_59;
 assign sub_860_43_n_56 = ~sub_860_43_n_55;
 assign sub_860_43_n_54 = ~sub_860_43_n_53;
 assign sub_860_43_n_52 = ~sub_860_43_n_51;
 assign sub_860_43_n_69 = (n_1178 | n_1293);
 assign sub_860_43_n_68 = ~(sub_860_43_n_50 & R_11_16_);
 assign sub_860_43_n_67 = ~(R_11_0_ & ~n_1351);
 assign sub_860_43_n_66 = ~(R_11_19_ | ~n_1213);
 assign sub_860_43_n_64 = ~(R_11_11_ | ~n_1027);
 assign sub_860_43_n_39 = ~(R_11_19_ & ~n_1213);
 assign sub_860_43_n_63 = ~(R_11_20_ | ~n_1367);
 assign sub_860_43_n_62 = ~(R_11_12_ | ~n_1260);
 assign sub_860_43_n_61 = ~(R_11_9_ | ~n_1346);
 assign sub_860_43_n_59 = ~(n_1341 | sub_860_43_n_48);
 assign sub_860_43_n_58 = ~(R_11_8_ | ~n_1163);
 assign sub_860_43_n_57 = ~(R_11_15_ | ~n_1137);
 assign sub_860_43_n_55 = ~(R_11_9_ & ~n_1346);
 assign sub_860_43_n_53 = ~(R_11_7_ | ~n_1218);
 assign sub_860_43_n_51 = ~(R_11_11_ & ~n_1027);
 assign sub_860_43_n_50 = ~n_1173;
 assign sub_860_43_n_49 = ~n_1168;
 assign sub_860_43_n_48 = ~R_11_3_;
 assign sub_860_43_n_47 = ~R_11_1_;
 assign sub_860_43_n_46 = ~R_11_16_;
 assign sub_860_43_n_38 = ~(n_1114 | ~R_11_2_);
 assign sub_860_43_n_37 = ~(n_1050 | ~R_11_4_);
 assign T_10_16_ = ~((sub_860_43_n_44 & ~sub_860_43_n_98) | (sub_860_43_n_157 & sub_860_43_n_98));
 assign sub_860_43_n_35 = ~(sub_860_43_n_150 & sub_860_43_n_129);
 assign sub_860_43_n_34 = ~(sub_860_43_n_118 & ~sub_860_43_n_117);
 assign sub_860_43_n_33 = ~(sub_860_43_n_140 | sub_860_43_n_106);
 assign sub_860_43_n_32 = ~(sub_860_43_n_35 & sub_860_43_n_102);
 assign sub_860_43_n_31 = ~(sub_860_43_n_145 & sub_860_43_n_94);
 assign sub_860_43_n_30 = ~(sub_860_43_n_71 | ~sub_860_43_n_4);
 assign sub_860_43_n_29 = (sub_860_43_n_60 & sub_860_43_n_5);
 assign sub_860_43_n_28 = ~(sub_860_43_n_37 | ~sub_860_43_n_11);
 assign sub_860_43_n_27 = ~(sub_860_43_n_14 & ~sub_860_43_n_83);
 assign sub_860_43_n_26 = ~(sub_860_43_n_83 | (sub_860_43_n_14 & sub_860_43_n_134));
 assign sub_860_43_n_25 = (sub_860_43_n_68 & sub_860_43_n_74);
 assign sub_860_43_n_24 = ~(sub_860_43_n_2 & ~sub_860_43_n_73);
 assign sub_860_43_n_23 = ~(sub_860_43_n_41 & (sub_860_43_n_72 | sub_860_43_n_167));
 assign sub_860_43_n_22 = ~(sub_860_43_n_62 | ~sub_860_43_n_3);
 assign sub_860_43_n_21 = ~(sub_860_43_n_82 | ~sub_860_43_n_6);
 assign sub_860_43_n_20 = ~(sub_860_43_n_39 & (sub_860_43_n_66 | sub_860_43_n_165));
 assign sub_860_43_n_19 = ~(sub_860_43_n_66 | ~sub_860_43_n_39);
 assign sub_860_43_n_18 = ~(sub_860_43_n_1 & ~sub_860_43_n_63);
 assign sub_860_43_n_17 = ~(sub_860_43_n_38 | ~sub_860_43_n_13);
 assign sub_860_43_n_16 = ~(sub_860_43_n_79 | ~sub_860_43_n_7);
 assign sub_860_43_n_15 = ~(sub_860_43_n_12 & ~sub_860_43_n_58);
 assign sub_860_43_n_14 = ~(sub_860_43_n_47 & n_1102);
 assign sub_860_43_n_13 = ~(n_1114 & ~R_11_2_);
 assign sub_860_43_n_12 = ~(R_11_8_ & ~n_1163);
 assign sub_860_43_n_11 = ~(n_1050 & ~R_11_4_);
 assign sub_860_43_n_10 = ~(R_11_18_ & ~n_1303);
 assign sub_860_43_n_9 = (R_11_6_ | sub_860_43_n_49);
 assign sub_860_43_n_8 = ~(R_11_7_ & ~n_1218);
 assign sub_860_43_n_7 = ~(n_1097 & ~R_11_5_);
 assign sub_860_43_n_6 = ~(R_11_14_ & ~n_1092);
 assign sub_860_43_n_5 = ~(sub_860_43_n_48 & n_1341);
 assign sub_860_43_n_4 = ~(R_11_10_ & ~n_1066);
 assign sub_860_43_n_3 = ~(R_11_12_ & ~n_1260);
 assign sub_860_43_n_2 = ~(R_11_13_ & ~n_1183);
 assign sub_860_43_n_1 = ~(R_11_20_ & ~n_1367);
 assign sub_860_43_n_0 = ~(n_1351 & ~R_11_0_);
 assign T_9_22_ = ((sub_890_40_n_31 & n_920) | ~(sub_890_40_n_31 | n_920));
 assign T_9_21_ = ((sub_890_40_n_192 & n_937) | ~(sub_890_40_n_192 | n_937));
 assign T_9_19_ = ~((sub_890_40_n_191 | n_919) & ~(sub_890_40_n_191 & n_919));
 assign T_9_15_ = ((sub_890_40_n_101 & ~sub_890_40_n_35) | (n_922 & sub_890_40_n_35));
 assign sub_890_40_n_192 = ~(n_927 & (~n_925 | n_962));
 assign sub_890_40_n_191 = ~(n_908 & (~n_959 | n_961));
 assign T_9_20_ = ~((sub_890_40_n_181 | sub_890_40_n_113) & ~(sub_890_40_n_181 & sub_890_40_n_113));
 assign T_9_18_ = ~((sub_890_40_n_183 | sub_890_40_n_98) & ~(sub_890_40_n_183 & sub_890_40_n_98));
 assign T_9_17_ = ~((n_914 | n_947) & ~(n_914 & n_947));
 assign T_9_14_ = ((n_916 & n_957) | ~(n_916 | n_957));
 assign T_9_13_ = ~((n_915 | n_946) & ~(n_915 & n_946));
 assign T_9_11_ = ~((n_932 | n_941) & ~(n_932 & n_941));
 assign sub_890_40_n_183 = ~n_961;
 assign sub_890_40_n_181 = ~n_962;
 assign sub_890_40_n_179 = ~(sub_890_40_n_158 & sub_890_40_n_172);
 assign sub_890_40_n_184 = ~(sub_890_40_n_71 & (~sub_890_40_n_85 | sub_890_40_n_169));
 assign sub_890_40_n_182 = ~(sub_890_40_n_173 | ~sub_890_40_n_128);
 assign sub_890_40_n_180 = ~(sub_890_40_n_145 | (~sub_890_40_n_138 & sub_890_40_n_170));
 assign T_9_10_ = ((sub_890_40_n_28 & sub_890_40_n_24) | ~(sub_890_40_n_28 | sub_890_40_n_24));
 assign T_9_12_ = ((sub_890_40_n_168 & sub_890_40_n_99) | ~(sub_890_40_n_168 | sub_890_40_n_99));
 assign T_9_7_ = ~((sub_890_40_n_171 | sub_890_40_n_14) & ~(sub_890_40_n_171 & sub_890_40_n_14));
 assign T_9_9_ = ((sub_890_40_n_167 & sub_890_40_n_17) | ~(sub_890_40_n_167 | sub_890_40_n_17));
 assign T_9_16_ = ((n_913 & n_939) | ~(n_913 | n_939));
 assign sub_890_40_n_173 = ~(sub_890_40_n_169 | ~sub_890_40_n_108);
 assign sub_890_40_n_172 = ~(sub_890_40_n_170 & ~sub_890_40_n_150);
 assign sub_890_40_n_171 = ~(sub_890_40_n_0 & (~sub_890_40_n_63 | sub_890_40_n_32));
 assign sub_890_40_n_169 = ~sub_890_40_n_170;
 assign sub_890_40_n_170 = ~(sub_890_40_n_163 & sub_890_40_n_152);
 assign sub_890_40_n_168 = ~(sub_890_40_n_164 & ~sub_890_40_n_144);
 assign sub_890_40_n_167 = ~(sub_890_40_n_13 & (~sub_890_40_n_59 | sub_890_40_n_38));
 assign T_9_6_ = ((sub_890_40_n_162 & sub_890_40_n_95) | ~(sub_890_40_n_162 | sub_890_40_n_95));
 assign T_9_5_ = ~((sub_890_40_n_21 | sub_890_40_n_20) & ~(sub_890_40_n_21 & sub_890_40_n_20));
 assign sub_890_40_n_164 = ~(sub_890_40_n_161 & ~sub_890_40_n_134);
 assign sub_890_40_n_163 = ~(sub_890_40_n_161 & sub_890_40_n_139);
 assign sub_890_40_n_162 = ~sub_890_40_n_32;
 assign sub_890_40_n_161 = ~(sub_890_40_n_143 & (sub_890_40_n_130 | sub_890_40_n_155));
 assign T_9_3_ = ((sub_890_40_n_23 & sub_890_40_n_16) | ~(sub_890_40_n_23 | sub_890_40_n_16));
 assign T_9_4_ = ((sub_890_40_n_157 & sub_890_40_n_18) | ~(sub_890_40_n_157 | sub_890_40_n_18));
 assign sub_890_40_n_158 = ~(sub_890_40_n_132 & (sub_890_40_n_149 | (sub_890_40_n_135 & sub_890_40_n_145)));
 assign sub_890_40_n_157 = ~sub_890_40_n_156;
 assign sub_890_40_n_156 = ~sub_890_40_n_155;
 assign sub_890_40_n_155 = ~(sub_890_40_n_129 | (sub_890_40_n_151 & sub_890_40_n_105));
 assign T_9_2_ = ~((sub_890_40_n_151 | sub_890_40_n_15) & ~(sub_890_40_n_151 & sub_890_40_n_15));
 assign sub_890_40_n_153 = ~(sub_890_40_n_151 & ~sub_890_40_n_50);
 assign sub_890_40_n_152 = ~(sub_890_40_n_146 | (sub_890_40_n_144 & sub_890_40_n_137));
 assign sub_890_40_n_151 = ~(sub_890_40_n_147 & sub_890_40_n_88);
 assign sub_890_40_n_150 = ~(sub_890_40_n_142 & sub_890_40_n_135);
 assign sub_890_40_n_149 = ~(sub_890_40_n_106 & (sub_890_40_n_126 | sub_890_40_n_117));
 assign T_9_1_ = ((sub_890_40_n_96 & n_1240) | ~(sub_890_40_n_96 | n_1240));
 assign sub_890_40_n_147 = ~(sub_890_40_n_141 | (n_1240 & R_10_0_));
 assign sub_890_40_n_146 = ~(sub_890_40_n_122 & (sub_890_40_n_125 | sub_890_40_n_115));
 assign sub_890_40_n_145 = ~(sub_890_40_n_124 & (~sub_890_40_n_104 | sub_890_40_n_128));
 assign sub_890_40_n_144 = ~(sub_890_40_n_140 & ~sub_890_40_n_123);
 assign sub_890_40_n_143 = ~(sub_890_40_n_121 | (sub_890_40_n_133 & sub_890_40_n_112));
 assign sub_890_40_n_142 = ~(sub_890_40_n_131 | sub_890_40_n_138);
 assign sub_890_40_n_141 = ~(n_1351 | ~n_1240);
 assign sub_890_40_n_140 = ~(sub_890_40_n_127 & sub_890_40_n_102);
 assign sub_890_40_n_139 = ~(sub_890_40_n_134 | sub_890_40_n_136);
 assign sub_890_40_n_137 = ~sub_890_40_n_136;
 assign sub_890_40_n_132 = ~sub_890_40_n_131;
 assign sub_890_40_n_130 = ~(sub_890_40_n_118 & sub_890_40_n_112);
 assign sub_890_40_n_129 = ~(sub_890_40_n_11 & (sub_890_40_n_43 | sub_890_40_n_51));
 assign sub_890_40_n_138 = ~(sub_890_40_n_104 & sub_890_40_n_108);
 assign sub_890_40_n_136 = ~(sub_890_40_n_110 & sub_890_40_n_114);
 assign sub_890_40_n_135 = ~(sub_890_40_n_116 | sub_890_40_n_117);
 assign sub_890_40_n_134 = ~(sub_890_40_n_97 & sub_890_40_n_102);
 assign sub_890_40_n_133 = ~(sub_890_40_n_2 & (sub_890_40_n_40 | sub_890_40_n_64));
 assign sub_890_40_n_131 = ~(sub_890_40_n_91 & sub_890_40_n_94);
 assign sub_890_40_n_124 = ~(sub_890_40_n_69 | (sub_890_40_n_65 & sub_890_40_n_77));
 assign sub_890_40_n_123 = ~(sub_890_40_n_87 & (sub_890_40_n_9 | sub_890_40_n_79));
 assign sub_890_40_n_122 = ~(sub_890_40_n_90 | (sub_890_40_n_53 & sub_890_40_n_81));
 assign sub_890_40_n_121 = ~(sub_890_40_n_3 & (sub_890_40_n_0 | sub_890_40_n_49));
 assign sub_890_40_n_128 = ~(sub_890_40_n_92 | ~sub_890_40_n_86);
 assign sub_890_40_n_127 = ~(sub_890_40_n_4 & (sub_890_40_n_13 | sub_890_40_n_52));
 assign sub_890_40_n_126 = ~(sub_890_40_n_107 | ~sub_890_40_n_68);
 assign sub_890_40_n_125 = ~(sub_890_40_n_12 | (sub_890_40_n_61 & sub_890_40_n_74));
 assign sub_890_40_n_115 = ~sub_890_40_n_114;
 assign sub_890_40_n_107 = ~(sub_890_40_n_66 | ~sub_890_40_n_57);
 assign sub_890_40_n_106 = ~(sub_890_40_n_6 & ~n_1293);
 assign sub_890_40_n_105 = ~(sub_890_40_n_50 | sub_890_40_n_51);
 assign sub_890_40_n_120 = ~(sub_890_40_n_5 & sub_890_40_n_73);
 assign sub_890_40_n_119 = ~(sub_890_40_n_86 & sub_890_40_n_67);
 assign sub_890_40_n_118 = ~(sub_890_40_n_78 | sub_890_40_n_64);
 assign sub_890_40_n_117 = ~(sub_890_40_n_10 & ~n_1293);
 assign sub_890_40_n_116 = ~(sub_890_40_n_8 & ~sub_890_40_n_56);
 assign sub_890_40_n_114 = ~(sub_890_40_n_72 | sub_890_40_n_80);
 assign sub_890_40_n_113 = ~(n_927 & n_925);
 assign sub_890_40_n_112 = ~(sub_890_40_n_62 | sub_890_40_n_49);
 assign sub_890_40_n_111 = ~(sub_890_40_n_68 & sub_890_40_n_57);
 assign sub_890_40_n_110 = ~(sub_890_40_n_54 | sub_890_40_n_60);
 assign sub_890_40_n_109 = ~(sub_890_40_n_1 & sub_890_40_n_77);
 assign sub_890_40_n_108 = ~(sub_890_40_n_84 | ~sub_890_40_n_67);
 assign sub_890_40_n_101 = ~n_922;
 assign sub_890_40_n_94 = ~(n_1298 | (n_1362 | (n_831 | n_1274)));
 assign T_9_0_ = ~(sub_890_40_n_70 & (~{in2[9]} | {in1[0]}));
 assign sub_890_40_n_92 = ~(sub_890_40_n_71 | ~sub_890_40_n_67);
 assign sub_890_40_n_91 = ~(n_1060 | (n_1372 | (n_1087 | n_1243)));
 assign sub_890_40_n_104 = ~(sub_890_40_n_82 | sub_890_40_n_76);
 assign sub_890_40_n_103 = ~(sub_890_40_n_13 & sub_890_40_n_59);
 assign sub_890_40_n_102 = ~(sub_890_40_n_41 | sub_890_40_n_79);
 assign sub_890_40_n_100 = ~(sub_890_40_n_89 & sub_890_40_n_81);
 assign sub_890_40_n_99 = ~(sub_890_40_n_75 & sub_890_40_n_55);
 assign sub_890_40_n_98 = ~(n_908 & n_959);
 assign sub_890_40_n_97 = ~(sub_890_40_n_58 | sub_890_40_n_52);
 assign sub_890_40_n_96 = ~(sub_890_40_n_88 & sub_890_40_n_7);
 assign sub_890_40_n_95 = ~(sub_890_40_n_0 & sub_890_40_n_63);
 assign sub_890_40_n_90 = ~sub_890_40_n_89;
 assign sub_890_40_n_85 = ~sub_890_40_n_84;
 assign sub_890_40_n_83 = ~sub_890_40_n_82;
 assign sub_890_40_n_81 = ~sub_890_40_n_80;
 assign sub_890_40_n_77 = ~sub_890_40_n_76;
 assign sub_890_40_n_75 = ~sub_890_40_n_74;
 assign sub_890_40_n_73 = ~sub_890_40_n_72;
 assign sub_890_40_n_89 = ~(sub_890_40_n_46 & R_10_14_);
 assign sub_890_40_n_88 = ~(R_10_0_ & ~n_1351);
 assign sub_890_40_n_87 = ~(R_10_10_ & ~n_1066);
 assign sub_890_40_n_86 = ~(sub_890_40_n_48 & sub_890_40_n_37);
 assign sub_890_40_n_84 = ~(R_10_15_ | ~n_1137);
 assign sub_890_40_n_82 = ~(R_10_17_ | ~n_1032);
 assign sub_890_40_n_80 = ~(R_10_14_ | ~n_1092);
 assign sub_890_40_n_43 = ~(R_10_1_ & ~n_1102);
 assign sub_890_40_n_79 = ~(R_10_10_ | ~n_1066);
 assign sub_890_40_n_78 = ~(R_10_3_ | ~n_1341);
 assign sub_890_40_n_76 = ~(R_10_18_ | ~n_1303);
 assign sub_890_40_n_74 = ~(n_1027 | sub_890_40_n_47);
 assign sub_890_40_n_72 = ~(R_10_13_ | ~n_1183);
 assign sub_890_40_n_71 = ~(sub_890_40_n_45 & R_10_15_);
 assign sub_890_40_n_70 = ~({in1[0]} & ~{in2[9]});
 assign sub_890_40_n_69 = ~sub_890_40_n_1;
 assign sub_890_40_n_65 = ~sub_890_40_n_42;
 assign sub_890_40_n_63 = ~sub_890_40_n_62;
 assign sub_890_40_n_61 = ~sub_890_40_n_60;
 assign sub_890_40_n_59 = ~sub_890_40_n_58;
 assign sub_890_40_n_57 = ~sub_890_40_n_56;
 assign sub_890_40_n_55 = ~sub_890_40_n_54;
 assign sub_890_40_n_53 = ~sub_890_40_n_5;
 assign sub_890_40_n_68 = ~(R_10_20_ & ~n_1367);
 assign sub_890_40_n_67 = ~(sub_890_40_n_36 & ~sub_890_40_n_48);
 assign sub_890_40_n_66 = ~(R_10_19_ & ~n_1213);
 assign sub_890_40_n_42 = ~(R_10_17_ & ~n_1032);
 assign sub_890_40_n_64 = ~(R_10_4_ | ~n_1050);
 assign sub_890_40_n_62 = ~(R_10_5_ | ~n_1097);
 assign sub_890_40_n_60 = ~(R_10_12_ | ~n_1260);
 assign sub_890_40_n_58 = ~(R_10_7_ | ~n_1218);
 assign sub_890_40_n_41 = ~(R_10_9_ | ~n_1346);
 assign sub_890_40_n_56 = ~(R_10_20_ | ~n_1367);
 assign sub_890_40_n_54 = ~(R_10_11_ | ~n_1027);
 assign sub_890_40_n_40 = ~(R_10_3_ & ~n_1341);
 assign sub_890_40_n_52 = ~(R_10_8_ | ~n_1163);
 assign sub_890_40_n_51 = ~(R_10_2_ | ~n_1114);
 assign sub_890_40_n_50 = ~(R_10_1_ | ~n_1102);
 assign sub_890_40_n_49 = ~(R_10_6_ | ~n_1168);
 assign sub_890_40_n_48 = ~n_1173;
 assign sub_890_40_n_47 = ~R_10_11_;
 assign sub_890_40_n_46 = ~n_1092;
 assign sub_890_40_n_45 = ~n_1137;
 assign T_9_32_ = ~n_909;
 assign sub_890_40_n_38 = ~sub_890_40_n_161;
 assign sub_890_40_n_37 = ~sub_890_40_n_36;
 assign sub_890_40_n_36 = ~R_10_16_;
 assign sub_890_40_n_35 = ~(n_956 & ~(n_958 & n_916));
 assign sub_890_40_n_34 = ~(sub_890_40_n_75 & ~(sub_890_40_n_55 & sub_890_40_n_168));
 assign sub_890_40_n_33 = ~(sub_890_40_n_30 & sub_890_40_n_125);
 assign sub_890_40_n_32 = ~(sub_890_40_n_133 | (sub_890_40_n_118 & sub_890_40_n_156));
 assign sub_890_40_n_31 = ~(n_928 & (n_963 | n_962));
 assign sub_890_40_n_30 = ~(sub_890_40_n_168 & sub_890_40_n_110);
 assign T_9_8_ = (sub_890_40_n_38 ^ sub_890_40_n_103);
 assign sub_890_40_n_28 = ~(sub_890_40_n_127 | (sub_890_40_n_97 & sub_890_40_n_161));
 assign sub_890_40_n_27 = ~(sub_890_40_n_61 & ~sub_890_40_n_12);
 assign sub_890_40_n_26 = ~(sub_890_40_n_10 & ~sub_890_40_n_6);
 assign sub_890_40_n_25 = (sub_890_40_n_71 & sub_890_40_n_85);
 assign sub_890_40_n_24 = ~(sub_890_40_n_41 | ~sub_890_40_n_9);
 assign sub_890_40_n_23 = ~(sub_890_40_n_153 & sub_890_40_n_43);
 assign sub_890_40_n_22 = ~(sub_890_40_n_87 & ~sub_890_40_n_79);
 assign sub_890_40_n_21 = ~(sub_890_40_n_40 & (sub_890_40_n_78 | sub_890_40_n_157));
 assign sub_890_40_n_20 = ~(sub_890_40_n_2 & ~sub_890_40_n_64);
 assign sub_890_40_n_19 = ~(sub_890_40_n_9 & (sub_890_40_n_41 | sub_890_40_n_28));
 assign sub_890_40_n_18 = ~(sub_890_40_n_78 | ~sub_890_40_n_40);
 assign sub_890_40_n_17 = ~(sub_890_40_n_4 & ~sub_890_40_n_52);
 assign sub_890_40_n_16 = ~(sub_890_40_n_11 & ~sub_890_40_n_51);
 assign sub_890_40_n_15 = ~(sub_890_40_n_43 & ~sub_890_40_n_50);
 assign sub_890_40_n_14 = ~(sub_890_40_n_3 & ~sub_890_40_n_49);
 assign sub_890_40_n_13 = ~(R_10_7_ & ~n_1218);
 assign sub_890_40_n_12 = ~(n_1260 | ~R_10_12_);
 assign sub_890_40_n_11 = ~(R_10_2_ & ~n_1114);
 assign sub_890_40_n_10 = ~(n_1178 & ~R_10_21_);
 assign sub_890_40_n_9 = ~(R_10_9_ & ~n_1346);
 assign sub_890_40_n_8 = ~(n_1213 & ~R_10_19_);
 assign sub_890_40_n_7 = ~(n_1351 & ~R_10_0_);
 assign sub_890_40_n_6 = ~(n_1178 | ~R_10_21_);
 assign sub_890_40_n_5 = ~(R_10_13_ & ~n_1183);
 assign sub_890_40_n_4 = ~(R_10_8_ & ~n_1163);
 assign sub_890_40_n_3 = ~(R_10_6_ & ~n_1168);
 assign sub_890_40_n_2 = ~(R_10_4_ & ~n_1050);
 assign sub_890_40_n_1 = ~(R_10_18_ & ~n_1303);
 assign sub_890_40_n_0 = ~(R_10_5_ & ~n_1097);
 assign T_8_23_ = ((sub_920_38_n_27 & sub_920_38_n_25) | ~(sub_920_38_n_27 | sub_920_38_n_25));
 assign T_8_21_ = ((sub_920_38_n_21 & ~sub_920_38_n_213) | (sub_920_38_n_115 & sub_920_38_n_213));
 assign T_8_19_ = ((sub_920_38_n_19 & ~sub_920_38_n_212) | (sub_920_38_n_33 & sub_920_38_n_212));
 assign T_8_15_ = ~((sub_920_38_n_215 | sub_920_38_n_28) & ~(sub_920_38_n_215 & sub_920_38_n_28));
 assign T_8_22_ = ((sub_920_38_n_200 & sub_920_38_n_32) | ~(sub_920_38_n_200 | sub_920_38_n_32));
 assign sub_920_38_n_213 = ~(sub_920_38_n_79 | (~sub_920_38_n_67 & sub_920_38_n_199));
 assign sub_920_38_n_215 = ~(sub_920_38_n_84 | (~sub_920_38_n_85 & sub_920_38_n_201));
 assign sub_920_38_n_212 = ~(sub_920_38_n_68 | (~sub_920_38_n_61 & sub_920_38_n_196));
 assign T_8_20_ = ((sub_920_38_n_199 & sub_920_38_n_22) | ~(sub_920_38_n_199 | sub_920_38_n_22));
 assign T_8_18_ = ((sub_920_38_n_196 & sub_920_38_n_20) | ~(sub_920_38_n_196 | sub_920_38_n_20));
 assign T_8_17_ = ((sub_920_38_n_197 & sub_920_38_n_30) | ~(sub_920_38_n_197 | sub_920_38_n_30));
 assign T_8_14_ = ~((sub_920_38_n_202 | sub_920_38_n_105) & ~(sub_920_38_n_202 & sub_920_38_n_105));
 assign T_8_13_ = ~((sub_920_38_n_204 | sub_920_38_n_36) & ~(sub_920_38_n_204 & sub_920_38_n_36));
 assign T_8_11_ = ~((sub_920_38_n_203 | sub_920_38_n_23) & ~(sub_920_38_n_203 & sub_920_38_n_23));
 assign T_8_32_ = ~sub_920_38_n_198;
 assign sub_920_38_n_202 = ~sub_920_38_n_201;
 assign sub_920_38_n_198 = ~(sub_920_38_n_190 & ~sub_920_38_n_173);
 assign sub_920_38_n_204 = ~(sub_920_38_n_75 | (~sub_920_38_n_82 & sub_920_38_n_184));
 assign sub_920_38_n_203 = ~(sub_920_38_n_6 | (~sub_920_38_n_91 & sub_920_38_n_38));
 assign sub_920_38_n_201 = ~(sub_920_38_n_134 & (~sub_920_38_n_114 | sub_920_38_n_39));
 assign sub_920_38_n_200 = ~(sub_920_38_n_129 | (sub_920_38_n_185 & sub_920_38_n_167));
 assign sub_920_38_n_199 = ~(sub_920_38_n_156 & (~sub_920_38_n_138 | sub_920_38_n_189));
 assign T_8_16_ = ((sub_920_38_n_189 & sub_920_38_n_110) | ~(sub_920_38_n_189 | sub_920_38_n_110));
 assign T_8_12_ = ((sub_920_38_n_39 & sub_920_38_n_106) | ~(sub_920_38_n_39 | sub_920_38_n_106));
 assign T_8_10_ = ~((sub_920_38_n_187 | sub_920_38_n_122) & ~(sub_920_38_n_187 & sub_920_38_n_122));
 assign T_8_9_ = ~((sub_920_38_n_186 | sub_920_38_n_24) & ~(sub_920_38_n_186 & sub_920_38_n_24));
 assign T_8_7_ = ~((sub_920_38_n_31 | sub_920_38_n_29) & ~(sub_920_38_n_31 & sub_920_38_n_29));
 assign sub_920_38_n_197 = ~(sub_920_38_n_92 | (~sub_920_38_n_60 & sub_920_38_n_188));
 assign sub_920_38_n_196 = ~(sub_920_38_n_131 & (~sub_920_38_n_111 | sub_920_38_n_189));
 assign sub_920_38_n_190 = ~(sub_920_38_n_188 & ~sub_920_38_n_162);
 assign sub_920_38_n_189 = ~sub_920_38_n_188;
 assign sub_920_38_n_188 = ~(sub_920_38_n_168 & sub_920_38_n_179);
 assign sub_920_38_n_187 = ~sub_920_38_n_38;
 assign sub_920_38_n_186 = ~(sub_920_38_n_41 | (~sub_920_38_n_66 & sub_920_38_n_178));
 assign sub_920_38_n_185 = ~(sub_920_38_n_179 & sub_920_38_n_40);
 assign sub_920_38_n_184 = ~sub_920_38_n_39;
 assign T_8_6_ = ~((sub_920_38_n_37 | sub_920_38_n_102) & ~(sub_920_38_n_37 & sub_920_38_n_102));
 assign T_8_5_ = ~((sub_920_38_n_176 | sub_920_38_n_34) & ~(sub_920_38_n_176 & sub_920_38_n_34));
 assign T_8_8_ = ((sub_920_38_n_178 & sub_920_38_n_121) | ~(sub_920_38_n_178 | sub_920_38_n_121));
 assign sub_920_38_n_180 = ~(sub_920_38_n_178 & ~sub_920_38_n_108);
 assign sub_920_38_n_179 = ~(sub_920_38_n_178 & ~sub_920_38_n_147);
 assign sub_920_38_n_178 = ~(sub_920_38_n_159 & (sub_920_38_n_42 | sub_920_38_n_136));
 assign sub_920_38_n_177 = ~(sub_920_38_n_140 & (~sub_920_38_n_123 | sub_920_38_n_42));
 assign sub_920_38_n_176 = ~(sub_920_38_n_88 | (~sub_920_38_n_89 & sub_920_38_n_171));
 assign T_8_4_ = ~((sub_920_38_n_172 | sub_920_38_n_116) & ~(sub_920_38_n_172 & sub_920_38_n_116));
 assign T_8_3_ = ~((sub_920_38_n_170 | sub_920_38_n_35) & ~(sub_920_38_n_170 & sub_920_38_n_35));
 assign sub_920_38_n_173 = ~(sub_920_38_n_142 | (sub_920_38_n_152 & (sub_920_38_n_154 | sub_920_38_n_143)));
 assign sub_920_38_n_172 = ~sub_920_38_n_171;
 assign sub_920_38_n_171 = ~sub_920_38_n_42;
 assign sub_920_38_n_42 = ~(sub_920_38_n_126 | (sub_920_38_n_165 & sub_920_38_n_164));
 assign sub_920_38_n_170 = ~(sub_920_38_n_80 | (~sub_920_38_n_73 & sub_920_38_n_166));
 assign T_8_2_ = ~((sub_920_38_n_166 | sub_920_38_n_26) & ~(sub_920_38_n_166 & sub_920_38_n_26));
 assign sub_920_38_n_168 = ~(sub_920_38_n_158 | (sub_920_38_n_153 & sub_920_38_n_145));
 assign sub_920_38_n_167 = ~(sub_920_38_n_118 | (~sub_920_38_n_138 & sub_920_38_n_156));
 assign sub_920_38_n_166 = ~(sub_920_38_n_150 & (sub_920_38_n_148 & sub_920_38_n_77));
 assign sub_920_38_n_165 = ~(sub_920_38_n_73 | ~sub_920_38_n_161);
 assign sub_920_38_n_164 = ~(sub_920_38_n_163 | sub_920_38_n_94);
 assign sub_920_38_n_163 = ~(sub_920_38_n_149 | R_9_0_);
 assign sub_920_38_n_162 = ~(sub_920_38_n_151 & sub_920_38_n_144);
 assign sub_920_38_n_161 = ~(sub_920_38_n_146 & (n_1352 & sub_920_38_n_150));
 assign T_8_1_ = ((sub_920_38_n_103 & n_1199) | ~(sub_920_38_n_103 | n_1199));
 assign sub_920_38_n_159 = ~(sub_920_38_n_135 | (sub_920_38_n_112 & sub_920_38_n_139));
 assign sub_920_38_n_158 = ~sub_920_38_n_157;
 assign sub_920_38_n_157 = ~(sub_920_38_n_124 | (sub_920_38_n_133 & sub_920_38_n_120));
 assign sub_920_38_n_156 = ~sub_920_38_n_155;
 assign sub_920_38_n_155 = ~sub_920_38_n_154;
 assign sub_920_38_n_154 = ~(sub_920_38_n_128 | (sub_920_38_n_130 & sub_920_38_n_107));
 assign sub_920_38_n_153 = ~(sub_920_38_n_125 & (sub_920_38_n_132 | sub_920_38_n_109));
 assign sub_920_38_n_152 = ~(sub_920_38_n_127 | (sub_920_38_n_129 & sub_920_38_n_104));
 assign sub_920_38_n_151 = ~(sub_920_38_n_142 | sub_920_38_n_137);
 assign sub_920_38_n_150 = ~sub_920_38_n_149;
 assign sub_920_38_n_149 = ~(sub_920_38_n_146 | n_1352);
 assign sub_920_38_n_148 = ~(R_9_0_ & ~sub_920_38_n_146);
 assign sub_920_38_n_147 = ~(sub_920_38_n_141 & sub_920_38_n_145);
 assign sub_920_38_n_146 = ~n_1199;
 assign sub_920_38_n_144 = ~sub_920_38_n_143;
 assign sub_920_38_n_140 = ~sub_920_38_n_139;
 assign sub_920_38_n_138 = ~sub_920_38_n_137;
 assign sub_920_38_n_136 = ~(sub_920_38_n_123 & sub_920_38_n_112);
 assign sub_920_38_n_135 = ~(sub_920_38_n_13 & (sub_920_38_n_64 | sub_920_38_n_90));
 assign sub_920_38_n_145 = ~(sub_920_38_n_113 | sub_920_38_n_119);
 assign sub_920_38_n_143 = ~(sub_920_38_n_117 & sub_920_38_n_104);
 assign sub_920_38_n_142 = ~(sub_920_38_n_99 & sub_920_38_n_100);
 assign sub_920_38_n_141 = ~(sub_920_38_n_109 | sub_920_38_n_108);
 assign sub_920_38_n_139 = ~(sub_920_38_n_18 & (sub_920_38_n_17 | sub_920_38_n_63));
 assign sub_920_38_n_137 = ~(sub_920_38_n_111 & sub_920_38_n_107);
 assign sub_920_38_n_134 = ~sub_920_38_n_133;
 assign sub_920_38_n_131 = ~sub_920_38_n_130;
 assign sub_920_38_n_128 = ~(sub_920_38_n_95 & (sub_920_38_n_11 | sub_920_38_n_58));
 assign sub_920_38_n_127 = ~(sub_920_38_n_1 & (sub_920_38_n_12 | sub_920_38_n_70));
 assign sub_920_38_n_126 = ~(sub_920_38_n_2 & (sub_920_38_n_4 | sub_920_38_n_94));
 assign sub_920_38_n_125 = ~(sub_920_38_n_97 | (sub_920_38_n_6 & sub_920_38_n_5));
 assign sub_920_38_n_124 = ~(sub_920_38_n_14 & (sub_920_38_n_83 | sub_920_38_n_87));
 assign sub_920_38_n_133 = ~(sub_920_38_n_98 & (sub_920_38_n_74 | sub_920_38_n_59));
 assign sub_920_38_n_132 = ~(sub_920_38_n_0 | (sub_920_38_n_41 & sub_920_38_n_10));
 assign sub_920_38_n_130 = ~(sub_920_38_n_8 & (sub_920_38_n_16 | sub_920_38_n_72));
 assign sub_920_38_n_129 = ~(sub_920_38_n_96 & (sub_920_38_n_78 | sub_920_38_n_62));
 assign sub_920_38_n_120 = ~sub_920_38_n_119;
 assign sub_920_38_n_118 = ~sub_920_38_n_117;
 assign sub_920_38_n_115 = ~sub_920_38_n_21;
 assign sub_920_38_n_114 = ~sub_920_38_n_113;
 assign sub_920_38_n_123 = ~(sub_920_38_n_89 | sub_920_38_n_63);
 assign sub_920_38_n_122 = ~(sub_920_38_n_6 | sub_920_38_n_91);
 assign sub_920_38_n_121 = ~(sub_920_38_n_69 & sub_920_38_n_9);
 assign sub_920_38_n_119 = ~(sub_920_38_n_86 & sub_920_38_n_3);
 assign sub_920_38_n_117 = ~(sub_920_38_n_67 | sub_920_38_n_62);
 assign sub_920_38_n_116 = ~(sub_920_38_n_88 | sub_920_38_n_89);
 assign sub_920_38_n_113 = ~(sub_920_38_n_81 & ~sub_920_38_n_56);
 assign sub_920_38_n_112 = ~(sub_920_38_n_93 | sub_920_38_n_90);
 assign sub_920_38_n_111 = ~(sub_920_38_n_60 | ~sub_920_38_n_71);
 assign T_8_0_ = ~(sub_920_38_n_57 & (~{in2[8]} | {in1[0]}));
 assign sub_920_38_n_100 = ~(n_1299 | (n_1363 | (n_832 | n_1275)));
 assign sub_920_38_n_99 = ~(n_1061 | (n_1373 | (n_1088 | n_1244)));
 assign sub_920_38_n_110 = ~(sub_920_38_n_92 | sub_920_38_n_60);
 assign sub_920_38_n_109 = ~(sub_920_38_n_15 & sub_920_38_n_5);
 assign sub_920_38_n_108 = ~(sub_920_38_n_9 & sub_920_38_n_10);
 assign sub_920_38_n_107 = ~(sub_920_38_n_61 | sub_920_38_n_58);
 assign sub_920_38_n_106 = ~(sub_920_38_n_75 | sub_920_38_n_82);
 assign sub_920_38_n_105 = ~(sub_920_38_n_84 | sub_920_38_n_85);
 assign sub_920_38_n_104 = ~(sub_920_38_n_76 | sub_920_38_n_70);
 assign sub_920_38_n_103 = ~(sub_920_38_n_77 & sub_920_38_n_7);
 assign sub_920_38_n_102 = ~(sub_920_38_n_65 | sub_920_38_n_93);
 assign sub_920_38_n_92 = ~sub_920_38_n_16;
 assign sub_920_38_n_91 = ~sub_920_38_n_15;
 assign sub_920_38_n_88 = ~sub_920_38_n_17;
 assign sub_920_38_n_87 = ~sub_920_38_n_86;
 assign sub_920_38_n_85 = ~sub_920_38_n_3;
 assign sub_920_38_n_84 = ~sub_920_38_n_83;
 assign sub_920_38_n_82 = ~sub_920_38_n_81;
 assign sub_920_38_n_80 = ~sub_920_38_n_4;
 assign sub_920_38_n_79 = ~sub_920_38_n_78;
 assign sub_920_38_n_98 = ~(sub_920_38_n_45 & R_9_12_);
 assign sub_920_38_n_97 = ~(n_1067 | sub_920_38_n_55);
 assign sub_920_38_n_96 = ~(R_9_20_ & ~n_1368);
 assign sub_920_38_n_95 = ~(R_9_18_ & ~n_1304);
 assign sub_920_38_n_94 = ~(R_9_2_ | ~n_1115);
 assign sub_920_38_n_93 = ~(R_9_5_ | ~n_1098);
 assign sub_920_38_n_90 = ~(R_9_6_ | ~n_1169);
 assign sub_920_38_n_89 = ~(R_9_3_ | ~n_1342);
 assign sub_920_38_n_86 = ~(sub_920_38_n_54 & ~sub_920_38_n_49);
 assign sub_920_38_n_83 = ~(sub_920_38_n_47 & ~n_1184);
 assign sub_920_38_n_81 = ~(sub_920_38_n_53 & ~sub_920_38_n_52);
 assign sub_920_38_n_78 = ~(R_9_19_ & ~n_1214);
 assign sub_920_38_n_75 = ~sub_920_38_n_74;
 assign sub_920_38_n_72 = ~sub_920_38_n_71;
 assign sub_920_38_n_69 = ~sub_920_38_n_41;
 assign sub_920_38_n_68 = ~sub_920_38_n_11;
 assign sub_920_38_n_66 = ~sub_920_38_n_9;
 assign sub_920_38_n_65 = ~sub_920_38_n_64;
 assign sub_920_38_n_77 = ~(sub_920_38_n_44 & R_9_0_);
 assign sub_920_38_n_76 = ~(R_9_21_ | ~n_1179);
 assign sub_920_38_n_74 = ~(sub_920_38_n_52 & R_9_11_);
 assign sub_920_38_n_73 = ~(R_9_1_ | ~n_1103);
 assign sub_920_38_n_71 = ~(sub_920_38_n_51 & ~sub_920_38_n_50);
 assign sub_920_38_n_70 = ~(R_9_22_ | ~n_1294);
 assign sub_920_38_n_41 = ~(n_1219 | sub_920_38_n_48);
 assign sub_920_38_n_67 = ~(R_9_19_ | ~n_1214);
 assign sub_920_38_n_64 = ~(R_9_5_ & ~n_1098);
 assign sub_920_38_n_63 = ~(R_9_4_ | ~n_1051);
 assign sub_920_38_n_62 = ~(R_9_20_ | ~n_1368);
 assign sub_920_38_n_61 = ~(R_9_17_ | ~n_1033);
 assign sub_920_38_n_60 = ~(R_9_15_ | ~n_1138);
 assign sub_920_38_n_56 = ~(R_9_12_ | ~n_1261);
 assign sub_920_38_n_59 = ~(R_9_12_ | ~n_1261);
 assign sub_920_38_n_58 = ~(R_9_18_ | ~n_1304);
 assign sub_920_38_n_57 = ~({in1[0]} & ~{in2[8]});
 assign sub_920_38_n_55 = ~R_9_10_;
 assign sub_920_38_n_54 = ~R_9_14_;
 assign sub_920_38_n_53 = ~R_9_11_;
 assign sub_920_38_n_52 = ~n_1028;
 assign sub_920_38_n_51 = ~R_9_16_;
 assign sub_920_38_n_50 = ~n_1174;
 assign sub_920_38_n_49 = ~n_1093;
 assign sub_920_38_n_48 = ~R_9_7_;
 assign sub_920_38_n_47 = ~sub_920_38_n_46;
 assign sub_920_38_n_46 = ~R_9_13_;
 assign sub_920_38_n_45 = ~n_1261;
 assign sub_920_38_n_44 = ~n_1352;
 assign sub_920_38_n_40 = ~(sub_920_38_n_155 | ~sub_920_38_n_168);
 assign sub_920_38_n_39 = ~(sub_920_38_n_153 | (sub_920_38_n_141 & sub_920_38_n_178));
 assign sub_920_38_n_38 = ~(sub_920_38_n_180 & sub_920_38_n_132);
 assign sub_920_38_n_37 = ~(sub_920_38_n_139 | (sub_920_38_n_123 & sub_920_38_n_171));
 assign sub_920_38_n_36 = ~(sub_920_38_n_59 | ~sub_920_38_n_98);
 assign sub_920_38_n_35 = ~(sub_920_38_n_94 | ~sub_920_38_n_2);
 assign sub_920_38_n_34 = ~(sub_920_38_n_63 | ~sub_920_38_n_18);
 assign sub_920_38_n_33 = ~(sub_920_38_n_58 | ~sub_920_38_n_95);
 assign sub_920_38_n_32 = ~(sub_920_38_n_76 | ~sub_920_38_n_12);
 assign sub_920_38_n_31 = ~(sub_920_38_n_65 | (~sub_920_38_n_93 & sub_920_38_n_177));
 assign sub_920_38_n_30 = ~(sub_920_38_n_72 | ~sub_920_38_n_8);
 assign sub_920_38_n_29 = ~(sub_920_38_n_90 | ~sub_920_38_n_13);
 assign sub_920_38_n_28 = ~(sub_920_38_n_87 | ~sub_920_38_n_14);
 assign sub_920_38_n_27 = ~(sub_920_38_n_12 & (sub_920_38_n_76 | sub_920_38_n_200));
 assign sub_920_38_n_26 = ~(sub_920_38_n_4 & ~sub_920_38_n_73);
 assign sub_920_38_n_25 = ~(sub_920_38_n_1 & ~sub_920_38_n_70);
 assign sub_920_38_n_24 = ~(sub_920_38_n_0 | ~sub_920_38_n_10);
 assign sub_920_38_n_23 = ~(sub_920_38_n_97 | ~sub_920_38_n_5);
 assign sub_920_38_n_22 = ~(sub_920_38_n_78 & ~sub_920_38_n_67);
 assign sub_920_38_n_21 = ~(sub_920_38_n_96 & ~sub_920_38_n_62);
 assign sub_920_38_n_20 = ~(sub_920_38_n_11 & ~sub_920_38_n_61);
 assign sub_920_38_n_19 = ~(sub_920_38_n_95 & ~sub_920_38_n_58);
 assign sub_920_38_n_18 = ~(R_9_4_ & ~n_1051);
 assign sub_920_38_n_17 = ~(R_9_3_ & ~n_1342);
 assign sub_920_38_n_16 = ~(R_9_15_ & ~n_1138);
 assign sub_920_38_n_15 = ~(n_1347 & ~R_9_9_);
 assign sub_920_38_n_14 = ~(sub_920_38_n_49 & ~sub_920_38_n_54);
 assign sub_920_38_n_13 = ~(R_9_6_ & ~n_1169);
 assign sub_920_38_n_12 = ~(R_9_21_ & ~n_1179);
 assign sub_920_38_n_11 = ~(R_9_17_ & ~n_1033);
 assign sub_920_38_n_10 = ~(n_1164 & ~R_9_8_);
 assign sub_920_38_n_9 = ~(sub_920_38_n_48 & n_1219);
 assign sub_920_38_n_8 = ~(sub_920_38_n_50 & ~sub_920_38_n_51);
 assign sub_920_38_n_7 = (R_9_0_ | sub_920_38_n_44);
 assign sub_920_38_n_6 = ~(n_1347 | ~R_9_9_);
 assign sub_920_38_n_5 = ~(sub_920_38_n_55 & n_1067);
 assign sub_920_38_n_4 = ~(R_9_1_ & ~n_1103);
 assign sub_920_38_n_3 = ~(sub_920_38_n_46 & n_1184);
 assign sub_920_38_n_2 = ~(R_9_2_ & ~n_1115);
 assign sub_920_38_n_1 = ~(R_9_22_ & ~n_1294);
 assign sub_920_38_n_0 = ~(n_1164 | ~R_9_8_);
 assign T_7_23_ = ((sub_950_37_n_201 & sub_950_37_n_37) | ~(sub_950_37_n_201 | sub_950_37_n_37));
 assign T_7_22_ = ((sub_950_37_n_203 & sub_950_37_n_112) | ~(sub_950_37_n_203 | sub_950_37_n_112));
 assign T_7_21_ = ((sub_950_37_n_26 & sub_950_37_n_103) | ~(sub_950_37_n_26 | sub_950_37_n_103));
 assign T_7_19_ = ((sub_950_37_n_202 & sub_950_37_n_19) | ~(sub_950_37_n_202 | sub_950_37_n_19));
 assign T_7_15_ = ((sub_950_37_n_25 & sub_950_37_n_30) | ~(sub_950_37_n_25 | sub_950_37_n_30));
 assign T_7_11_ = ((sub_950_37_n_189 & sub_950_37_n_32) | ~(sub_950_37_n_189 | sub_950_37_n_32));
 assign sub_950_37_n_203 = ~(sub_950_37_n_193 & ~sub_950_37_n_120);
 assign sub_950_37_n_202 = ~(sub_950_37_n_191 & ~sub_950_37_n_71);
 assign sub_950_37_n_201 = ~(sub_950_37_n_70 & (sub_950_37_n_143 | (sub_950_37_n_176 & sub_950_37_n_145)));
 assign T_7_24_ = ((sub_950_37_n_188 & sub_950_37_n_45) | ~(sub_950_37_n_188 | sub_950_37_n_45));
 assign T_7_20_ = ((sub_950_37_n_187 & sub_950_37_n_40) | ~(sub_950_37_n_187 | sub_950_37_n_40));
 assign T_7_17_ = ((sub_950_37_n_185 & sub_950_37_n_46) | ~(sub_950_37_n_185 | sub_950_37_n_46));
 assign T_7_18_ = ((sub_950_37_n_53 & sub_950_37_n_35) | ~(sub_950_37_n_53 | sub_950_37_n_35));
 assign T_7_14_ = ((sub_950_37_n_184 & sub_950_37_n_31) | ~(sub_950_37_n_184 | sub_950_37_n_31));
 assign T_7_13_ = ((sub_950_37_n_39 & sub_950_37_n_27) | ~(sub_950_37_n_39 | sub_950_37_n_27));
 assign sub_950_37_n_193 = ~(sub_950_37_n_187 & ~sub_950_37_n_110);
 assign sub_950_37_n_192 = ~(sub_950_37_n_187 & ~sub_950_37_n_86);
 assign sub_950_37_n_191 = ~(sub_950_37_n_53 & ~sub_950_37_n_82);
 assign sub_950_37_n_190 = ~(sub_950_37_n_184 & ~sub_950_37_n_79);
 assign T_7_32_ = ~(sub_950_37_n_174 | sub_950_37_n_157);
 assign sub_950_37_n_189 = ~(sub_950_37_n_18 & ~sub_950_37_n_89);
 assign sub_950_37_n_188 = ~(sub_950_37_n_177 & ~sub_950_37_n_150);
 assign sub_950_37_n_187 = ~(sub_950_37_n_176 & ~sub_950_37_n_140);
 assign T_7_16_ = ~((sub_950_37_n_173 | sub_950_37_n_24) & ~(sub_950_37_n_173 & sub_950_37_n_24));
 assign T_7_7_ = ((sub_950_37_n_20 & sub_950_37_n_17) | ~(sub_950_37_n_20 | sub_950_37_n_17));
 assign T_7_12_ = ((sub_950_37_n_169 & sub_950_37_n_34) | ~(sub_950_37_n_169 | sub_950_37_n_34));
 assign T_7_10_ = ((sub_950_37_n_52 & sub_950_37_n_42) | ~(sub_950_37_n_52 | sub_950_37_n_42));
 assign T_7_9_ = ((sub_950_37_n_170 & sub_950_37_n_33) | ~(sub_950_37_n_170 | sub_950_37_n_33));
 assign sub_950_37_n_185 = ~(sub_950_37_n_29 & ~sub_950_37_n_7);
 assign sub_950_37_n_184 = ~(sub_950_37_n_49 & ~sub_950_37_n_124);
 assign sub_950_37_n_178 = ~(sub_950_37_n_169 & ~sub_950_37_n_81);
 assign sub_950_37_n_177 = ~(sub_950_37_n_173 & ~sub_950_37_n_136);
 assign sub_950_37_n_176 = ~(sub_950_37_n_172 & ~sub_950_37_n_134);
 assign sub_950_37_n_175 = ~(sub_950_37_n_173 & ~sub_950_37_n_111);
 assign sub_950_37_n_174 = ~(sub_950_37_n_171 | ~sub_950_37_n_144);
 assign sub_950_37_n_173 = ~sub_950_37_n_171;
 assign sub_950_37_n_172 = ~sub_950_37_n_171;
 assign sub_950_37_n_171 = ~(sub_950_37_n_151 | (sub_950_37_n_162 & sub_950_37_n_135));
 assign sub_950_37_n_170 = ~(sub_950_37_n_164 & ~sub_950_37_n_93);
 assign sub_950_37_n_169 = ~(sub_950_37_n_163 & ~sub_950_37_n_139);
 assign T_7_6_ = ~((sub_950_37_n_161 | sub_950_37_n_22) & ~(sub_950_37_n_161 & sub_950_37_n_22));
 assign T_7_5_ = ~((sub_950_37_n_28 | sub_950_37_n_38) & ~(sub_950_37_n_28 & sub_950_37_n_38));
 assign T_7_8_ = ((sub_950_37_n_162 & sub_950_37_n_44) | ~(sub_950_37_n_162 | sub_950_37_n_44));
 assign sub_950_37_n_165 = ~(sub_950_37_n_161 & ~sub_950_37_n_73);
 assign sub_950_37_n_164 = ~(sub_950_37_n_162 & ~sub_950_37_n_3);
 assign sub_950_37_n_163 = ~(sub_950_37_n_162 & ~sub_950_37_n_133);
 assign sub_950_37_n_162 = ~(sub_950_37_n_142 & sub_950_37_n_158);
 assign sub_950_37_n_161 = ~(sub_950_37_n_48 & ~sub_950_37_n_123);
 assign T_7_4_ = ~((sub_950_37_n_155 | sub_950_37_n_41) & ~(sub_950_37_n_155 & sub_950_37_n_41));
 assign sub_950_37_n_159 = ~(sub_950_37_n_155 & ~sub_950_37_n_88);
 assign sub_950_37_n_158 = ~(sub_950_37_n_155 & ~sub_950_37_n_128);
 assign sub_950_37_n_157 = ~(sub_950_37_n_156 & ~sub_950_37_n_54);
 assign sub_950_37_n_156 = ~(sub_950_37_n_150 & ~sub_950_37_n_138);
 assign sub_950_37_n_155 = ~(sub_950_37_n_152 & sub_950_37_n_116);
 assign T_7_2_ = ~((sub_950_37_n_149 | sub_950_37_n_36) & ~(sub_950_37_n_149 & sub_950_37_n_36));
 assign sub_950_37_n_153 = ~(sub_950_37_n_149 & ~sub_950_37_n_83);
 assign sub_950_37_n_152 = ~(sub_950_37_n_149 & sub_950_37_n_107);
 assign sub_950_37_n_151 = ~(sub_950_37_n_146 & sub_950_37_n_141);
 assign sub_950_37_n_150 = ~(sub_950_37_n_147 & sub_950_37_n_56);
 assign sub_950_37_n_149 = ((n_1150 & R_8_0_) | ((R_8_0_ & sub_950_37_n_65) | (sub_950_37_n_65 & n_1150)));
 assign T_7_1_ = (R_8_0_ ^ (sub_950_37_n_65 ^ n_1150));
 assign sub_950_37_n_147 = ~(sub_950_37_n_140 & ~sub_950_37_n_130);
 assign sub_950_37_n_146 = ~(sub_950_37_n_139 & ~sub_950_37_n_129);
 assign sub_950_37_n_145 = ~(sub_950_37_n_140 | ~sub_950_37_n_119);
 assign sub_950_37_n_144 = ~(sub_950_37_n_136 | ~sub_950_37_n_137);
 assign sub_950_37_n_143 = ~(sub_950_37_n_92 & (sub_950_37_n_120 | sub_950_37_n_59));
 assign sub_950_37_n_142 = ~(sub_950_37_n_127 | (sub_950_37_n_123 & sub_950_37_n_104));
 assign sub_950_37_n_141 = ~(sub_950_37_n_126 | (sub_950_37_n_124 & sub_950_37_n_113));
 assign sub_950_37_n_140 = ~(sub_950_37_n_55 & (~sub_950_37_n_100 | sub_950_37_n_122));
 assign sub_950_37_n_139 = ~(sub_950_37_n_118 & (sub_950_37_n_121 | sub_950_37_n_101));
 assign sub_950_37_n_138 = ~sub_950_37_n_137;
 assign sub_950_37_n_137 = ~(sub_950_37_n_94 | ~sub_950_37_n_132);
 assign sub_950_37_n_136 = ~(sub_950_37_n_47 & sub_950_37_n_131);
 assign sub_950_37_n_135 = ~(sub_950_37_n_133 | sub_950_37_n_129);
 assign sub_950_37_n_134 = ~sub_950_37_n_47;
 assign sub_950_37_n_131 = ~sub_950_37_n_130;
 assign sub_950_37_n_128 = ~(sub_950_37_n_105 & sub_950_37_n_104);
 assign sub_950_37_n_127 = ~(sub_950_37_n_13 & (sub_950_37_n_1 | sub_950_37_n_69));
 assign sub_950_37_n_126 = ~(sub_950_37_n_12 & (sub_950_37_n_74 | sub_950_37_n_77));
 assign sub_950_37_n_133 = ~(sub_950_37_n_23 & sub_950_37_n_102);
 assign sub_950_37_n_132 = ~(n_1088 | (n_1244 | (n_1275 | sub_950_37_n_98)));
 assign sub_950_37_n_130 = ~(sub_950_37_n_59 & sub_950_37_n_114);
 assign sub_950_37_n_129 = ~(sub_950_37_n_106 & sub_950_37_n_113);
 assign sub_950_37_n_125 = ~sub_950_37_n_117;
 assign sub_950_37_n_120 = ~sub_950_37_n_119;
 assign sub_950_37_n_118 = ~(sub_950_37_n_80 | (sub_950_37_n_89 & sub_950_37_n_8));
 assign sub_950_37_n_117 = ~(sub_950_37_n_97 & (sub_950_37_n_70 | sub_950_37_n_84));
 assign sub_950_37_n_116 = ~(sub_950_37_n_108 | ~sub_950_37_n_95);
 assign sub_950_37_n_124 = ~(sub_950_37_n_2 & (sub_950_37_n_58 | sub_950_37_n_76));
 assign sub_950_37_n_123 = ~(sub_950_37_n_6 & (sub_950_37_n_57 | sub_950_37_n_85));
 assign sub_950_37_n_122 = ~(sub_950_37_n_9 | (~sub_950_37_n_87 & sub_950_37_n_7));
 assign sub_950_37_n_121 = ~(sub_950_37_n_16 | (sub_950_37_n_93 & sub_950_37_n_15));
 assign sub_950_37_n_119 = ~(sub_950_37_n_109 | ~sub_950_37_n_96);
 assign sub_950_37_n_115 = ~sub_950_37_n_114;
 assign sub_950_37_n_110 = ~sub_950_37_n_59;
 assign sub_950_37_n_109 = ~(sub_950_37_n_75 | ~sub_950_37_n_78);
 assign sub_950_37_n_108 = ~(sub_950_37_n_0 | sub_950_37_n_90);
 assign sub_950_37_n_107 = ~(sub_950_37_n_83 | sub_950_37_n_90);
 assign sub_950_37_n_114 = ~(sub_950_37_n_91 | sub_950_37_n_84);
 assign sub_950_37_n_113 = ~(sub_950_37_n_79 | sub_950_37_n_77);
 assign sub_950_37_n_112 = ~(sub_950_37_n_70 & sub_950_37_n_92);
 assign sub_950_37_n_111 = ~(sub_950_37_n_10 & ~sub_950_37_n_87);
 assign sub_950_37_n_59 = ~(sub_950_37_n_86 | ~sub_950_37_n_78);
 assign sub_950_37_n_102 = ~sub_950_37_n_101;
 assign T_7_0_ = ~(sub_950_37_n_68 & (~{in2[7]} | {in1[0]}));
 assign sub_950_37_n_98 = (n_1373 | (n_1299 | (n_1363 | n_832)));
 assign sub_950_37_n_106 = ~(sub_950_37_n_81 | sub_950_37_n_76);
 assign sub_950_37_n_105 = ~(sub_950_37_n_88 | sub_950_37_n_85);
 assign sub_950_37_n_104 = ~(sub_950_37_n_73 | sub_950_37_n_69);
 assign sub_950_37_n_103 = ~(sub_950_37_n_96 & sub_950_37_n_78);
 assign sub_950_37_n_101 = ~(sub_950_37_n_4 & sub_950_37_n_8);
 assign sub_950_37_n_100 = ~(sub_950_37_n_82 | sub_950_37_n_72);
 assign sub_950_37_n_92 = ~sub_950_37_n_91;
 assign sub_950_37_n_97 = ~(R_8_22_ & ~n_1294);
 assign sub_950_37_n_96 = ~(sub_950_37_n_64 & ~n_1368);
 assign sub_950_37_n_95 = ~(R_8_2_ & ~n_1115);
 assign sub_950_37_n_94 = ~(R_8_23_ | ~n_1061);
 assign sub_950_37_n_93 = ~(n_1219 | sub_950_37_n_62);
 assign sub_950_37_n_91 = ~(R_8_21_ | ~n_1179);
 assign sub_950_37_n_90 = ~(R_8_2_ | ~n_1115);
 assign sub_950_37_n_89 = ~(n_1347 | sub_950_37_n_67);
 assign sub_950_37_n_88 = ~(R_8_3_ | ~n_1342);
 assign sub_950_37_n_87 = ~(R_8_16_ | ~n_1174);
 assign sub_950_37_n_86 = ~(R_8_19_ | ~n_1214);
 assign sub_950_37_n_58 = ~(R_8_11_ & ~n_1028);
 assign sub_950_37_n_85 = ~(R_8_4_ | ~n_1051);
 assign sub_950_37_n_84 = ~(R_8_22_ | ~n_1294);
 assign sub_950_37_n_83 = ~(R_8_1_ | ~n_1103);
 assign sub_950_37_n_82 = ~(R_8_17_ | ~n_1033);
 assign sub_950_37_n_81 = ~(R_8_11_ | ~n_1028);
 assign sub_950_37_n_71 = ~sub_950_37_n_11;
 assign sub_950_37_n_80 = ~(n_1067 | sub_950_37_n_66);
 assign sub_950_37_n_79 = ~(R_8_13_ | ~n_1184);
 assign sub_950_37_n_78 = ~(sub_950_37_n_63 & ~sub_950_37_n_61);
 assign sub_950_37_n_77 = ~(R_8_14_ | ~n_1093);
 assign sub_950_37_n_57 = ~(R_8_3_ & ~n_1342);
 assign sub_950_37_n_76 = ~(R_8_12_ | ~n_1261);
 assign sub_950_37_n_75 = ~(R_8_19_ & ~n_1214);
 assign sub_950_37_n_74 = ~(R_8_13_ & ~n_1184);
 assign sub_950_37_n_73 = ~(R_8_5_ | ~n_1098);
 assign sub_950_37_n_72 = ~(R_8_18_ | ~n_1304);
 assign sub_950_37_n_70 = ~(R_8_21_ & ~n_1179);
 assign sub_950_37_n_69 = ~(R_8_6_ | ~n_1169);
 assign sub_950_37_n_68 = ~({in1[0]} & ~{in2[7]});
 assign sub_950_37_n_67 = ~R_8_9_;
 assign sub_950_37_n_66 = ~R_8_10_;
 assign sub_950_37_n_65 = ~n_1352;
 assign sub_950_37_n_64 = ~sub_950_37_n_63;
 assign sub_950_37_n_63 = ~R_8_20_;
 assign sub_950_37_n_62 = ~R_8_7_;
 assign sub_950_37_n_61 = ~n_1368;
 assign sub_950_37_n_56 = (sub_950_37_n_125 & (sub_950_37_n_119 | sub_950_37_n_115));
 assign sub_950_37_n_55 = (sub_950_37_n_5 & (sub_950_37_n_11 | sub_950_37_n_72));
 assign sub_950_37_n_54 = ~(sub_950_37_n_14 | ~sub_950_37_n_132);
 assign sub_950_37_n_53 = ~(sub_950_37_n_175 & sub_950_37_n_122);
 assign sub_950_37_n_52 = ~(sub_950_37_n_51 & sub_950_37_n_121);
 assign sub_950_37_n_51 = ~(sub_950_37_n_162 & sub_950_37_n_23);
 assign T_7_3_ = ~(sub_950_37_n_21 ^ sub_950_37_n_43);
 assign sub_950_37_n_49 = ~(sub_950_37_n_169 & sub_950_37_n_106);
 assign sub_950_37_n_48 = ~(sub_950_37_n_155 & sub_950_37_n_105);
 assign sub_950_37_n_47 = ~(sub_950_37_n_111 | ~sub_950_37_n_100);
 assign sub_950_37_n_46 = (sub_950_37_n_9 | sub_950_37_n_87);
 assign sub_950_37_n_45 = ~(sub_950_37_n_14 & ~sub_950_37_n_94);
 assign sub_950_37_n_44 = (sub_950_37_n_93 | sub_950_37_n_3);
 assign sub_950_37_n_43 = ~(sub_950_37_n_95 & ~sub_950_37_n_90);
 assign sub_950_37_n_42 = ~(sub_950_37_n_4 & ~sub_950_37_n_89);
 assign sub_950_37_n_41 = ~(sub_950_37_n_57 & ~sub_950_37_n_88);
 assign sub_950_37_n_40 = ~(sub_950_37_n_75 & ~sub_950_37_n_86);
 assign sub_950_37_n_39 = ~(sub_950_37_n_178 & sub_950_37_n_58);
 assign sub_950_37_n_38 = ~(sub_950_37_n_6 & ~sub_950_37_n_85);
 assign sub_950_37_n_37 = ~(sub_950_37_n_97 & ~sub_950_37_n_84);
 assign sub_950_37_n_36 = ~(sub_950_37_n_0 & ~sub_950_37_n_83);
 assign sub_950_37_n_35 = ~(sub_950_37_n_11 & ~sub_950_37_n_82);
 assign sub_950_37_n_34 = ~(sub_950_37_n_58 & ~sub_950_37_n_81);
 assign sub_950_37_n_33 = ~(sub_950_37_n_15 & ~sub_950_37_n_16);
 assign sub_950_37_n_32 = ~(sub_950_37_n_8 & ~sub_950_37_n_80);
 assign sub_950_37_n_31 = ~(sub_950_37_n_74 & ~sub_950_37_n_79);
 assign sub_950_37_n_30 = ~(sub_950_37_n_12 & ~sub_950_37_n_77);
 assign sub_950_37_n_29 = ~(sub_950_37_n_173 & sub_950_37_n_10);
 assign sub_950_37_n_28 = ~(sub_950_37_n_159 & sub_950_37_n_57);
 assign sub_950_37_n_27 = ~(sub_950_37_n_2 & ~sub_950_37_n_76);
 assign sub_950_37_n_26 = ~(sub_950_37_n_192 & sub_950_37_n_75);
 assign sub_950_37_n_25 = ~(sub_950_37_n_190 & sub_950_37_n_74);
 assign sub_950_37_n_24 = ~(sub_950_37_n_10 & ~sub_950_37_n_7);
 assign sub_950_37_n_23 = ~(sub_950_37_n_3 | ~sub_950_37_n_15);
 assign sub_950_37_n_22 = ~(sub_950_37_n_1 & ~sub_950_37_n_73);
 assign sub_950_37_n_21 = ~(sub_950_37_n_153 & sub_950_37_n_0);
 assign sub_950_37_n_20 = ~(sub_950_37_n_165 & sub_950_37_n_1);
 assign sub_950_37_n_19 = ~(sub_950_37_n_5 & ~sub_950_37_n_72);
 assign sub_950_37_n_18 = ~(sub_950_37_n_52 & sub_950_37_n_4);
 assign sub_950_37_n_17 = ~(sub_950_37_n_13 & ~sub_950_37_n_69);
 assign sub_950_37_n_16 = ~(n_1164 | ~R_8_8_);
 assign sub_950_37_n_15 = ~(n_1164 & ~R_8_8_);
 assign sub_950_37_n_14 = ~(R_8_23_ & ~n_1061);
 assign sub_950_37_n_13 = ~(R_8_6_ & ~n_1169);
 assign sub_950_37_n_12 = ~(R_8_14_ & ~n_1093);
 assign sub_950_37_n_11 = ~(R_8_17_ & ~n_1033);
 assign sub_950_37_n_10 = ~(n_1138 & ~R_8_15_);
 assign sub_950_37_n_9 = ~(n_1174 | ~R_8_16_);
 assign sub_950_37_n_8 = ~(sub_950_37_n_66 & n_1067);
 assign sub_950_37_n_7 = ~(n_1138 | ~R_8_15_);
 assign sub_950_37_n_6 = ~(R_8_4_ & ~n_1051);
 assign sub_950_37_n_5 = ~(R_8_18_ & ~n_1304);
 assign sub_950_37_n_4 = ~(sub_950_37_n_67 & n_1347);
 assign sub_950_37_n_3 = (sub_950_37_n_62 & n_1219);
 assign sub_950_37_n_2 = ~(R_8_12_ & ~n_1261);
 assign sub_950_37_n_1 = ~(R_8_5_ & ~n_1098);
 assign sub_950_37_n_0 = ~(R_8_1_ & ~n_1103);
 assign T_6_25_ = ((sub_980_36_n_224 & sub_980_36_n_23) | ~(sub_980_36_n_224 | sub_980_36_n_23));
 assign T_6_23_ = ((sub_980_36_n_227 & sub_980_36_n_118) | ~(sub_980_36_n_227 | sub_980_36_n_118));
 assign T_6_21_ = ((sub_980_36_n_226 & sub_980_36_n_24) | ~(sub_980_36_n_226 | sub_980_36_n_24));
 assign T_6_19_ = ((sub_980_36_n_225 & sub_980_36_n_27) | ~(sub_980_36_n_225 | sub_980_36_n_27));
 assign T_6_15_ = ((sub_980_36_n_20 & sub_980_36_n_31) | ~(sub_980_36_n_20 | sub_980_36_n_31));
 assign T_6_14_ = ((sub_980_36_n_208 & sub_980_36_n_139) | ~(sub_980_36_n_208 | sub_980_36_n_139));
 assign sub_980_36_n_227 = ~(sub_980_36_n_44 & (sub_980_36_n_212 | sub_980_36_n_78));
 assign sub_980_36_n_226 = ~(sub_980_36_n_80 | (sub_980_36_n_38 & sub_980_36_n_43));
 assign sub_980_36_n_225 = ~(sub_980_36_n_98 | (~sub_980_36_n_93 & sub_980_36_n_211));
 assign sub_980_36_n_224 = ~(sub_980_36_n_103 | (sub_980_36_n_213 & sub_980_36_n_111));
 assign T_6_17_ = ((sub_980_36_n_209 & sub_980_36_n_28) | ~(sub_980_36_n_209 | sub_980_36_n_28));
 assign T_6_11_ = ((sub_980_36_n_215 & sub_980_36_n_29) | ~(sub_980_36_n_215 | sub_980_36_n_29));
 assign T_6_24_ = ((sub_980_36_n_213 & sub_980_36_n_123) | ~(sub_980_36_n_213 | sub_980_36_n_123));
 assign T_6_22_ = ((sub_980_36_n_212 & sub_980_36_n_127) | ~(sub_980_36_n_212 | sub_980_36_n_127));
 assign T_6_20_ = ((sub_980_36_n_48 & sub_980_36_n_17) | ~(sub_980_36_n_48 | sub_980_36_n_17));
 assign T_6_18_ = ((sub_980_36_n_211 & sub_980_36_n_122) | ~(sub_980_36_n_211 | sub_980_36_n_122));
 assign T_6_13_ = ((sub_980_36_n_214 & sub_980_36_n_30) | ~(sub_980_36_n_214 | sub_980_36_n_30));
 assign sub_980_36_n_48 = ~sub_980_36_n_38;
 assign T_6_32_ = ~(sub_980_36_n_197 | sub_980_36_n_182);
 assign sub_980_36_n_215 = ~(sub_980_36_n_101 | (~sub_980_36_n_109 & sub_980_36_n_196));
 assign sub_980_36_n_214 = ~(sub_980_36_n_74 | (~sub_980_36_n_72 & sub_980_36_n_37));
 assign sub_980_36_n_213 = ~(sub_980_36_n_201 & ~sub_980_36_n_176);
 assign sub_980_36_n_212 = ~(sub_980_36_n_35 | (~sub_980_36_n_161 & sub_980_36_n_194));
 assign sub_980_36_n_211 = ~(sub_980_36_n_199 & ~sub_980_36_n_154);
 assign sub_980_36_n_208 = ~sub_980_36_n_207;
 assign T_6_16_ = ~((sub_980_36_n_194 | sub_980_36_n_136) & ~(sub_980_36_n_194 & sub_980_36_n_136));
 assign T_6_7_ = ((sub_980_36_n_195 & sub_980_36_n_18) | ~(sub_980_36_n_195 | sub_980_36_n_18));
 assign T_6_12_ = ~((sub_980_36_n_37 | sub_980_36_n_21) & ~(sub_980_36_n_37 & sub_980_36_n_21));
 assign T_6_10_ = ~((sub_980_36_n_196 | sub_980_36_n_26) & ~(sub_980_36_n_196 & sub_980_36_n_26));
 assign T_6_9_ = ((sub_980_36_n_40 & sub_980_36_n_33) | ~(sub_980_36_n_40 | sub_980_36_n_33));
 assign sub_980_36_n_209 = ~(sub_980_36_n_95 | (~sub_980_36_n_96 & sub_980_36_n_194));
 assign sub_980_36_n_207 = ~(sub_980_36_n_198 & ~sub_980_36_n_149);
 assign sub_980_36_n_201 = ~(sub_980_36_n_194 & ~sub_980_36_n_163);
 assign sub_980_36_n_200 = ~(sub_980_36_n_194 & ~sub_980_36_n_153);
 assign sub_980_36_n_199 = ~(sub_980_36_n_194 & ~sub_980_36_n_119);
 assign sub_980_36_n_198 = ~(sub_980_36_n_37 & ~sub_980_36_n_126);
 assign sub_980_36_n_197 = ~(sub_980_36_n_193 | ~sub_980_36_n_174);
 assign sub_980_36_n_196 = ~(sub_980_36_n_147 & (~sub_980_36_n_134 | sub_980_36_n_47));
 assign sub_980_36_n_195 = ~(sub_980_36_n_69 | (~sub_980_36_n_81 & sub_980_36_n_34));
 assign sub_980_36_n_194 = ~sub_980_36_n_193;
 assign sub_980_36_n_193 = ~(sub_980_36_n_188 | sub_980_36_n_177);
 assign T_6_6_ = ((sub_980_36_n_185 & sub_980_36_n_133) | ~(sub_980_36_n_185 | sub_980_36_n_133));
 assign T_6_5_ = ((sub_980_36_n_39 & sub_980_36_n_25) | ~(sub_980_36_n_39 | sub_980_36_n_25));
 assign T_6_8_ = ((sub_980_36_n_47 & sub_980_36_n_135) | ~(sub_980_36_n_47 | sub_980_36_n_135));
 assign sub_980_36_n_189 = ~(sub_980_36_n_187 & ~sub_980_36_n_156);
 assign sub_980_36_n_188 = ~(sub_980_36_n_186 | ~sub_980_36_n_164);
 assign sub_980_36_n_47 = ~sub_980_36_n_187;
 assign sub_980_36_n_187 = ~sub_980_36_n_186;
 assign sub_980_36_n_186 = ~(sub_980_36_n_171 | (sub_980_36_n_179 & sub_980_36_n_151));
 assign sub_980_36_n_185 = ~sub_980_36_n_34;
 assign T_6_4_ = ((sub_980_36_n_46 & sub_980_36_n_121) | ~(sub_980_36_n_46 | sub_980_36_n_121));
 assign T_6_3_ = ((sub_980_36_n_180 & sub_980_36_n_19) | ~(sub_980_36_n_180 | sub_980_36_n_19));
 assign sub_980_36_n_182 = ~(sub_980_36_n_181 & ~sub_980_36_n_160);
 assign sub_980_36_n_181 = ~(sub_980_36_n_176 & ~sub_980_36_n_173);
 assign sub_980_36_n_180 = ~(sub_980_36_n_76 | (~sub_980_36_n_89 & sub_980_36_n_175));
 assign sub_980_36_n_46 = ~sub_980_36_n_179;
 assign sub_980_36_n_179 = ~(sub_980_36_n_142 & (sub_980_36_n_166 | sub_980_36_n_128));
 assign T_6_2_ = ~((sub_980_36_n_175 | sub_980_36_n_22) & ~(sub_980_36_n_175 & sub_980_36_n_22));
 assign sub_980_36_n_177 = ~(sub_980_36_n_170 & (sub_980_36_n_168 | sub_980_36_n_159));
 assign sub_980_36_n_176 = ~(sub_980_36_n_167 & (sub_980_36_n_158 | sub_980_36_n_169));
 assign sub_980_36_n_175 = ~sub_980_36_n_166;
 assign sub_980_36_n_174 = ~(sub_980_36_n_163 | ~sub_980_36_n_172);
 assign sub_980_36_n_173 = ~sub_980_36_n_172;
 assign sub_980_36_n_172 = ~(sub_980_36_n_155 | (sub_980_36_n_92 | sub_980_36_n_110));
 assign sub_980_36_n_171 = ~(sub_980_36_n_150 & (sub_980_36_n_137 | sub_980_36_n_148));
 assign sub_980_36_n_170 = ~(sub_980_36_n_143 | (sub_980_36_n_149 & sub_980_36_n_130));
 assign sub_980_36_n_169 = ~(sub_980_36_n_141 | (~sub_980_36_n_138 & sub_980_36_n_154));
 assign sub_980_36_n_168 = ~(sub_980_36_n_144 | (sub_980_36_n_146 & sub_980_36_n_120));
 assign sub_980_36_n_167 = ~(sub_980_36_n_140 | (sub_980_36_n_145 & sub_980_36_n_132));
 assign sub_980_36_n_166 = ~(sub_980_36_n_162 | ~sub_980_36_n_15);
 assign T_6_1_ = ((sub_980_36_n_32 & n_1228) | ~(sub_980_36_n_32 | n_1228));
 assign sub_980_36_n_164 = ~(sub_980_36_n_156 | sub_980_36_n_159);
 assign sub_980_36_n_163 = ~(sub_980_36_n_152 & sub_980_36_n_157);
 assign sub_980_36_n_162 = ~(sub_980_36_n_115 | ~n_1228);
 assign sub_980_36_n_161 = ~(sub_980_36_n_152 & ~sub_980_36_n_129);
 assign sub_980_36_n_160 = ~(sub_980_36_n_155 | (sub_980_36_n_6 & (sub_980_36_n_102 | sub_980_36_n_92)));
 assign sub_980_36_n_158 = ~sub_980_36_n_157;
 assign sub_980_36_n_153 = ~sub_980_36_n_152;
 assign sub_980_36_n_151 = ~(sub_980_36_n_124 | sub_980_36_n_137);
 assign sub_980_36_n_150 = ~(sub_980_36_n_90 | (sub_980_36_n_69 & sub_980_36_n_5));
 assign sub_980_36_n_159 = ~(sub_980_36_n_125 & sub_980_36_n_130);
 assign sub_980_36_n_157 = ~(sub_980_36_n_129 | sub_980_36_n_131);
 assign sub_980_36_n_156 = ~(sub_980_36_n_134 & sub_980_36_n_120);
 assign sub_980_36_n_155 = (n_832 | (n_1275 | sub_980_36_n_116));
 assign sub_980_36_n_154 = ~(sub_980_36_n_112 & (sub_980_36_n_94 | sub_980_36_n_99));
 assign sub_980_36_n_152 = ~(sub_980_36_n_138 | sub_980_36_n_119);
 assign sub_980_36_n_147 = ~sub_980_36_n_146;
 assign sub_980_36_n_144 = ~(sub_980_36_n_14 & (sub_980_36_n_8 | sub_980_36_n_73));
 assign sub_980_36_n_143 = ~(sub_980_36_n_1 & (sub_980_36_n_3 | sub_980_36_n_86));
 assign sub_980_36_n_142 = ~(sub_980_36_n_41 | (sub_980_36_n_4 & sub_980_36_n_76));
 assign sub_980_36_n_141 = ~(sub_980_36_n_12 & (sub_980_36_n_9 | sub_980_36_n_84));
 assign sub_980_36_n_140 = ~(sub_980_36_n_113 & (sub_980_36_n_44 | sub_980_36_n_104));
 assign sub_980_36_n_149 = ~(sub_980_36_n_10 & (sub_980_36_n_45 | sub_980_36_n_75));
 assign sub_980_36_n_148 = ~(sub_980_36_n_114 | (sub_980_36_n_42 & sub_980_36_n_100));
 assign sub_980_36_n_146 = ~(sub_980_36_n_0 & (sub_980_36_n_11 | sub_980_36_n_107));
 assign sub_980_36_n_145 = ~(sub_980_36_n_2 & (sub_980_36_n_79 | sub_980_36_n_87));
 assign sub_980_36_n_132 = ~sub_980_36_n_131;
 assign sub_980_36_n_128 = ~(sub_980_36_n_88 & sub_980_36_n_4);
 assign sub_980_36_n_139 = ~(sub_980_36_n_85 | sub_980_36_n_70);
 assign sub_980_36_n_138 = ~(sub_980_36_n_13 & sub_980_36_n_83);
 assign sub_980_36_n_137 = ~(sub_980_36_n_7 & sub_980_36_n_5);
 assign sub_980_36_n_136 = ~(sub_980_36_n_94 & sub_980_36_n_97);
 assign sub_980_36_n_135 = ~(sub_980_36_n_82 | sub_980_36_n_108);
 assign sub_980_36_n_134 = ~(sub_980_36_n_108 | sub_980_36_n_107);
 assign sub_980_36_n_133 = ~(sub_980_36_n_69 | sub_980_36_n_81);
 assign sub_980_36_n_131 = ~(sub_980_36_n_105 & sub_980_36_n_77);
 assign sub_980_36_n_130 = ~(sub_980_36_n_70 | sub_980_36_n_86);
 assign sub_980_36_n_129 = ~(sub_980_36_n_43 & ~sub_980_36_n_87);
 assign sub_980_36_n_126 = ~sub_980_36_n_125;
 assign T_6_0_ = ~(sub_980_36_n_68 & (~{in2[6]} | {in1[0]}));
 assign sub_980_36_n_116 = (n_1088 | (n_1244 | (n_1299 | n_1363)));
 assign sub_980_36_n_127 = ~(sub_980_36_n_71 | sub_980_36_n_78);
 assign sub_980_36_n_125 = ~(sub_980_36_n_72 | sub_980_36_n_75);
 assign sub_980_36_n_124 = ~(sub_980_36_n_16 & sub_980_36_n_100);
 assign sub_980_36_n_123 = ~(sub_980_36_n_102 & sub_980_36_n_111);
 assign sub_980_36_n_122 = ~(sub_980_36_n_9 & sub_980_36_n_13);
 assign sub_980_36_n_121 = ~(sub_980_36_n_42 | sub_980_36_n_106);
 assign sub_980_36_n_120 = ~(sub_980_36_n_109 | sub_980_36_n_73);
 assign sub_980_36_n_119 = ~(sub_980_36_n_97 & ~sub_980_36_n_99);
 assign sub_980_36_n_118 = ~(sub_980_36_n_113 & sub_980_36_n_105);
 assign sub_980_36_n_114 = ~sub_980_36_n_91;
 assign sub_980_36_n_111 = ~sub_980_36_n_110;
 assign sub_980_36_n_106 = ~sub_980_36_n_16;
 assign sub_980_36_n_104 = ~sub_980_36_n_105;
 assign sub_980_36_n_103 = ~sub_980_36_n_102;
 assign sub_980_36_n_101 = ~sub_980_36_n_8;
 assign sub_980_36_n_98 = ~sub_980_36_n_9;
 assign sub_980_36_n_96 = ~sub_980_36_n_97;
 assign sub_980_36_n_95 = ~sub_980_36_n_94;
 assign sub_980_36_n_93 = ~sub_980_36_n_13;
 assign sub_980_36_n_115 = ~(R_7_0_ | ~n_1352);
 assign sub_980_36_n_91 = ~(sub_980_36_n_63 & R_7_4_);
 assign sub_980_36_n_113 = ~(sub_980_36_n_66 & R_7_22_);
 assign sub_980_36_n_112 = ~(R_7_16_ & ~n_1174);
 assign sub_980_36_n_110 = ~(R_7_23_ | ~n_1061);
 assign sub_980_36_n_109 = ~(R_7_9_ | ~n_1347);
 assign sub_980_36_n_108 = ~(R_7_7_ | ~n_1219);
 assign sub_980_36_n_107 = ~(R_7_8_ | ~n_1164);
 assign sub_980_36_n_105 = ~(sub_980_36_n_56 & ~sub_980_36_n_66);
 assign sub_980_36_n_102 = ~(R_7_23_ & ~n_1061);
 assign sub_980_36_n_100 = ~(sub_980_36_n_57 & ~sub_980_36_n_63);
 assign sub_980_36_n_99 = ~(R_7_16_ | ~n_1174);
 assign sub_980_36_n_97 = ~(sub_980_36_n_65 & ~sub_980_36_n_51);
 assign sub_980_36_n_94 = ~(R_7_15_ & ~n_1138);
 assign sub_980_36_n_92 = ~(R_7_24_ | ~n_1373);
 assign sub_980_36_n_89 = ~sub_980_36_n_88;
 assign sub_980_36_n_85 = ~sub_980_36_n_3;
 assign sub_980_36_n_84 = ~sub_980_36_n_83;
 assign sub_980_36_n_82 = ~sub_980_36_n_11;
 assign sub_980_36_n_81 = ~sub_980_36_n_7;
 assign sub_980_36_n_80 = ~sub_980_36_n_79;
 assign sub_980_36_n_78 = ~sub_980_36_n_77;
 assign sub_980_36_n_74 = ~sub_980_36_n_45;
 assign sub_980_36_n_71 = ~sub_980_36_n_44;
 assign sub_980_36_n_90 = ~(n_1169 | sub_980_36_n_61);
 assign sub_980_36_n_88 = ~(sub_980_36_n_59 & ~sub_980_36_n_67);
 assign sub_980_36_n_87 = ~(R_7_20_ | ~n_1368);
 assign sub_980_36_n_86 = ~(R_7_14_ | ~n_1093);
 assign sub_980_36_n_83 = ~(sub_980_36_n_64 & ~sub_980_36_n_58);
 assign sub_980_36_n_79 = ~(R_7_19_ & ~n_1214);
 assign sub_980_36_n_77 = ~(sub_980_36_n_53 & ~sub_980_36_n_50);
 assign sub_980_36_n_76 = ~(n_1103 | sub_980_36_n_59);
 assign sub_980_36_n_75 = ~(R_7_12_ | ~n_1261);
 assign sub_980_36_n_45 = ~(R_7_11_ & ~n_1028);
 assign sub_980_36_n_73 = ~(R_7_10_ | ~n_1067);
 assign sub_980_36_n_72 = ~(R_7_11_ | ~n_1028);
 assign sub_980_36_n_44 = ~(sub_980_36_n_50 & sub_980_36_n_54);
 assign sub_980_36_n_70 = ~(R_7_13_ | ~n_1184);
 assign sub_980_36_n_69 = ~(n_1098 | sub_980_36_n_55);
 assign sub_980_36_n_43 = ~(sub_980_36_n_62 & ~sub_980_36_n_52);
 assign sub_980_36_n_68 = ~({in1[0]} & ~{in2[6]});
 assign sub_980_36_n_67 = ~n_1103;
 assign sub_980_36_n_66 = ~n_1294;
 assign sub_980_36_n_65 = ~R_7_15_;
 assign sub_980_36_n_64 = ~R_7_18_;
 assign sub_980_36_n_63 = ~n_1051;
 assign sub_980_36_n_62 = ~R_7_19_;
 assign sub_980_36_n_61 = ~R_7_6_;
 assign sub_980_36_n_60 = ~R_7_17_;
 assign sub_980_36_n_59 = ~R_7_1_;
 assign sub_980_36_n_58 = ~n_1304;
 assign sub_980_36_n_57 = ~R_7_4_;
 assign sub_980_36_n_56 = ~R_7_22_;
 assign sub_980_36_n_55 = ~R_7_5_;
 assign sub_980_36_n_54 = ~sub_980_36_n_53;
 assign sub_980_36_n_53 = ~R_7_21_;
 assign sub_980_36_n_52 = ~n_1214;
 assign sub_980_36_n_51 = ~n_1138;
 assign sub_980_36_n_50 = ~n_1179;
 assign sub_980_36_n_42 = ~(n_1342 | ~R_7_3_);
 assign sub_980_36_n_41 = ~(n_1115 | ~R_7_2_);
 assign sub_980_36_n_40 = ~(sub_980_36_n_82 | (~sub_980_36_n_108 & ~sub_980_36_n_47));
 assign sub_980_36_n_39 = ~(sub_980_36_n_42 | (~sub_980_36_n_106 & ~sub_980_36_n_46));
 assign sub_980_36_n_38 = ~(sub_980_36_n_200 & sub_980_36_n_169);
 assign sub_980_36_n_37 = ~(sub_980_36_n_189 & sub_980_36_n_168);
 assign sub_980_36_n_35 = ~sub_980_36_n_36;
 assign sub_980_36_n_36 = ~(sub_980_36_n_145 | (~sub_980_36_n_129 & ~sub_980_36_n_169));
 assign sub_980_36_n_34 = ~(sub_980_36_n_148 & (sub_980_36_n_124 | sub_980_36_n_46));
 assign sub_980_36_n_33 = ~(sub_980_36_n_107 | ~sub_980_36_n_0);
 assign sub_980_36_n_32 = ~(sub_980_36_n_15 & ~sub_980_36_n_115);
 assign sub_980_36_n_31 = ~(sub_980_36_n_86 | ~sub_980_36_n_1);
 assign sub_980_36_n_30 = ~(sub_980_36_n_75 | ~sub_980_36_n_10);
 assign sub_980_36_n_29 = ~(sub_980_36_n_73 | ~sub_980_36_n_14);
 assign sub_980_36_n_28 = ~(sub_980_36_n_99 | ~sub_980_36_n_112);
 assign sub_980_36_n_27 = ~(sub_980_36_n_84 | ~sub_980_36_n_12);
 assign sub_980_36_n_26 = ~(sub_980_36_n_8 & ~sub_980_36_n_109);
 assign sub_980_36_n_25 = ~(sub_980_36_n_114 | ~sub_980_36_n_100);
 assign sub_980_36_n_24 = ~(sub_980_36_n_87 | ~sub_980_36_n_2);
 assign sub_980_36_n_23 = ~(sub_980_36_n_92 | ~sub_980_36_n_6);
 assign sub_980_36_n_22 = (sub_980_36_n_76 | sub_980_36_n_89);
 assign sub_980_36_n_21 = ~(sub_980_36_n_45 & ~sub_980_36_n_72);
 assign sub_980_36_n_20 = ~(sub_980_36_n_85 | (~sub_980_36_n_70 & sub_980_36_n_207));
 assign sub_980_36_n_19 = ~(sub_980_36_n_41 | ~sub_980_36_n_4);
 assign sub_980_36_n_18 = ~(sub_980_36_n_90 | ~sub_980_36_n_5);
 assign sub_980_36_n_17 = ~(sub_980_36_n_80 | ~sub_980_36_n_43);
 assign sub_980_36_n_16 = ~(n_1342 & ~R_7_3_);
 assign sub_980_36_n_15 = ~(R_7_0_ & ~n_1352);
 assign sub_980_36_n_14 = ~(R_7_10_ & ~n_1067);
 assign sub_980_36_n_13 = ~(sub_980_36_n_60 & n_1033);
 assign sub_980_36_n_12 = ~(sub_980_36_n_58 & ~sub_980_36_n_64);
 assign sub_980_36_n_11 = ~(R_7_7_ & ~n_1219);
 assign sub_980_36_n_10 = ~(R_7_12_ & ~n_1261);
 assign sub_980_36_n_9 = (sub_980_36_n_60 | n_1033);
 assign sub_980_36_n_8 = ~(R_7_9_ & ~n_1347);
 assign sub_980_36_n_7 = ~(sub_980_36_n_55 & n_1098);
 assign sub_980_36_n_6 = ~(R_7_24_ & ~n_1373);
 assign sub_980_36_n_5 = ~(sub_980_36_n_61 & n_1169);
 assign sub_980_36_n_4 = ~(n_1115 & ~R_7_2_);
 assign sub_980_36_n_3 = ~(R_7_13_ & ~n_1184);
 assign sub_980_36_n_2 = ~(R_7_20_ & ~n_1368);
 assign sub_980_36_n_1 = ~(R_7_14_ & ~n_1093);
 assign sub_980_36_n_0 = ~(R_7_8_ & ~n_1164);
 assign T_5_26_ = ((sub_1010_35_n_234 & sub_1010_35_n_136) | ~(sub_1010_35_n_234 | sub_1010_35_n_136));
 assign T_5_15_ = ((sub_1010_35_n_35 & sub_1010_35_n_15) | ~(sub_1010_35_n_35 | sub_1010_35_n_15));
 assign T_5_25_ = ((sub_1010_35_n_233 & sub_1010_35_n_107) | ~(sub_1010_35_n_233 | sub_1010_35_n_107));
 assign T_5_21_ = ((sub_1010_35_n_232 & sub_1010_35_n_17) | ~(sub_1010_35_n_232 | sub_1010_35_n_17));
 assign T_5_19_ = ((sub_1010_35_n_231 & sub_1010_35_n_113) | ~(sub_1010_35_n_231 | sub_1010_35_n_113));
 assign T_5_23_ = ((sub_1010_35_n_21 & sub_1010_35_n_16) | ~(sub_1010_35_n_21 | sub_1010_35_n_16));
 assign T_5_14_ = ~((sub_1010_35_n_221 | sub_1010_35_n_140) & ~(sub_1010_35_n_221 & sub_1010_35_n_140));
 assign sub_1010_35_n_234 = ~(sub_1010_35_n_147 & (~sub_1010_35_n_111 | sub_1010_35_n_219));
 assign sub_1010_35_n_233 = ~(sub_1010_35_n_59 & (~sub_1010_35_n_38 | sub_1010_35_n_219));
 assign sub_1010_35_n_232 = ~(sub_1010_35_n_64 & (~sub_1010_35_n_92 | sub_1010_35_n_211));
 assign sub_1010_35_n_231 = ~(sub_1010_35_n_42 & (~sub_1010_35_n_72 | sub_1010_35_n_210));
 assign T_5_13_ = ((sub_1010_35_n_139 & ~sub_1010_35_n_34) | (sub_1010_35_n_20 & sub_1010_35_n_34));
 assign T_5_11_ = ~((sub_1010_35_n_25 | sub_1010_35_n_28) & ~(sub_1010_35_n_25 & sub_1010_35_n_28));
 assign T_5_24_ = ((sub_1010_35_n_220 & sub_1010_35_n_121) | ~(sub_1010_35_n_220 | sub_1010_35_n_121));
 assign T_5_20_ = ((sub_1010_35_n_217 & sub_1010_35_n_115) | ~(sub_1010_35_n_217 | sub_1010_35_n_115));
 assign T_5_18_ = ((sub_1010_35_n_32 & sub_1010_35_n_109) | ~(sub_1010_35_n_32 | sub_1010_35_n_109));
 assign T_5_17_ = ((sub_1010_35_n_222 & sub_1010_35_n_130) | ~(sub_1010_35_n_222 | sub_1010_35_n_130));
 assign T_5_22_ = ((sub_1010_35_n_47 & sub_1010_35_n_116) | ~(sub_1010_35_n_47 | sub_1010_35_n_116));
 assign sub_1010_35_n_219 = ~sub_1010_35_n_220;
 assign T_5_32_ = ~(sub_1010_35_n_207 | sub_1010_35_n_189);
 assign sub_1010_35_n_222 = ~(sub_1010_35_n_85 & (~sub_1010_35_n_70 | sub_1010_35_n_202));
 assign sub_1010_35_n_221 = ~(sub_1010_35_n_209 & ~sub_1010_35_n_150);
 assign sub_1010_35_n_220 = ~(sub_1010_35_n_208 & ~sub_1010_35_n_183);
 assign T_5_16_ = ((sub_1010_35_n_201 & sub_1010_35_n_127) | ~(sub_1010_35_n_201 | sub_1010_35_n_127));
 assign T_5_7_ = ~((sub_1010_35_n_203 | sub_1010_35_n_134) & ~(sub_1010_35_n_203 & sub_1010_35_n_134));
 assign T_5_12_ = ~((sub_1010_35_n_33 | sub_1010_35_n_137) & ~(sub_1010_35_n_33 & sub_1010_35_n_137));
 assign T_5_10_ = ((sub_1010_35_n_205 & sub_1010_35_n_19) | ~(sub_1010_35_n_205 | sub_1010_35_n_19));
 assign T_5_9_ = ~((sub_1010_35_n_204 | sub_1010_35_n_27) & ~(sub_1010_35_n_204 & sub_1010_35_n_27));
 assign sub_1010_35_n_211 = ~(sub_1010_35_n_167 | (~sub_1010_35_n_157 & sub_1010_35_n_201));
 assign sub_1010_35_n_217 = ~(sub_1010_35_n_168 & (~sub_1010_35_n_44 | sub_1010_35_n_202));
 assign sub_1010_35_n_210 = ~(sub_1010_35_n_152 | (~sub_1010_35_n_18 & sub_1010_35_n_201));
 assign sub_1010_35_n_209 = ~(sub_1010_35_n_33 & ~sub_1010_35_n_120);
 assign sub_1010_35_n_208 = ~(sub_1010_35_n_201 & ~sub_1010_35_n_164);
 assign sub_1010_35_n_207 = ~(sub_1010_35_n_202 | ~sub_1010_35_n_177);
 assign sub_1010_35_n_47 = ~sub_1010_35_n_206;
 assign sub_1010_35_n_206 = ~(sub_1010_35_n_197 | ~sub_1010_35_n_179);
 assign sub_1010_35_n_205 = ~(sub_1010_35_n_160 | (~sub_1010_35_n_142 & sub_1010_35_n_46));
 assign sub_1010_35_n_204 = ~(sub_1010_35_n_6 & (~sub_1010_35_n_97 | sub_1010_35_n_45));
 assign sub_1010_35_n_203 = ~(sub_1010_35_n_37 & (~sub_1010_35_n_3 | sub_1010_35_n_194));
 assign sub_1010_35_n_201 = ~sub_1010_35_n_202;
 assign sub_1010_35_n_202 = ~(sub_1010_35_n_196 | sub_1010_35_n_181);
 assign T_5_6_ = ~((sub_1010_35_n_30 | sub_1010_35_n_133) & ~(sub_1010_35_n_30 & sub_1010_35_n_133));
 assign T_5_5_ = ((sub_1010_35_n_192 & sub_1010_35_n_132) | ~(sub_1010_35_n_192 | sub_1010_35_n_132));
 assign T_5_8_ = ~((sub_1010_35_n_46 | sub_1010_35_n_135) & ~(sub_1010_35_n_46 & sub_1010_35_n_135));
 assign sub_1010_35_n_197 = ~(sub_1010_35_n_188 & (sub_1010_35_n_45 | sub_1010_35_n_176));
 assign sub_1010_35_n_196 = ~(sub_1010_35_n_45 | ~sub_1010_35_n_165);
 assign sub_1010_35_n_195 = ~(sub_1010_35_n_193 & ~sub_1010_35_n_159);
 assign sub_1010_35_n_194 = ~(sub_1010_35_n_149 | (~sub_1010_35_n_114 & sub_1010_35_n_187));
 assign sub_1010_35_n_46 = ~sub_1010_35_n_45;
 assign sub_1010_35_n_193 = ~sub_1010_35_n_45;
 assign sub_1010_35_n_45 = ~(sub_1010_35_n_171 | (sub_1010_35_n_187 & sub_1010_35_n_156));
 assign sub_1010_35_n_192 = ~(sub_1010_35_n_40 & (~sub_1010_35_n_5 | sub_1010_35_n_186));
 assign T_5_4_ = ((sub_1010_35_n_186 & sub_1010_35_n_23) | ~(sub_1010_35_n_186 | sub_1010_35_n_23));
 assign T_5_3_ = ((sub_1010_35_n_24 & sub_1010_35_n_22) | ~(sub_1010_35_n_24 | sub_1010_35_n_22));
 assign sub_1010_35_n_189 = ((sub_1010_35_n_175 & sub_1010_35_n_105) | ~(sub_1010_35_n_182 | sub_1010_35_n_163));
 assign sub_1010_35_n_188 = ~(sub_1010_35_n_181 & sub_1010_35_n_31);
 assign sub_1010_35_n_186 = ~sub_1010_35_n_187;
 assign sub_1010_35_n_187 = ~(sub_1010_35_n_180 & sub_1010_35_n_144);
 assign T_5_2_ = ~((sub_1010_35_n_178 | sub_1010_35_n_26) & ~(sub_1010_35_n_178 & sub_1010_35_n_26));
 assign sub_1010_35_n_184 = ~(sub_1010_35_n_178 & ~sub_1010_35_n_90);
 assign sub_1010_35_n_183 = ~sub_1010_35_n_182;
 assign sub_1010_35_n_182 = ~(sub_1010_35_n_172 | (sub_1010_35_n_161 & sub_1010_35_n_167));
 assign sub_1010_35_n_181 = ~(sub_1010_35_n_170 & (sub_1010_35_n_169 | sub_1010_35_n_158));
 assign sub_1010_35_n_180 = ~(sub_1010_35_n_178 & sub_1010_35_n_123);
 assign sub_1010_35_n_179 = ~(sub_1010_35_n_154 | (~sub_1010_35_n_126 & sub_1010_35_n_167));
 assign sub_1010_35_n_178 = ~(sub_1010_35_n_174 & sub_1010_35_n_78);
 assign sub_1010_35_n_177 = ~(sub_1010_35_n_164 | ~sub_1010_35_n_162);
 assign sub_1010_35_n_176 = ~(sub_1010_35_n_165 & sub_1010_35_n_31);
 assign sub_1010_35_n_175 = ~(sub_1010_35_n_29 & (sub_1010_35_n_147 | sub_1010_35_n_131));
 assign sub_1010_35_n_174 = ~(sub_1010_35_n_166 | (n_1042 & R_6_0_));
 assign T_5_1_ = ((sub_1010_35_n_108 & n_1042) | ~(sub_1010_35_n_108 | n_1042));
 assign sub_1010_35_n_172 = ~(sub_1010_35_n_36 & (sub_1010_35_n_153 | sub_1010_35_n_128));
 assign sub_1010_35_n_171 = ~(sub_1010_35_n_155 & (sub_1010_35_n_148 | sub_1010_35_n_138));
 assign sub_1010_35_n_170 = ~(sub_1010_35_n_143 | (sub_1010_35_n_150 & sub_1010_35_n_112));
 assign sub_1010_35_n_169 = ~(sub_1010_35_n_145 | (sub_1010_35_n_160 & sub_1010_35_n_129));
 assign sub_1010_35_n_168 = ~sub_1010_35_n_167;
 assign sub_1010_35_n_167 = ~(sub_1010_35_n_146 & (~sub_1010_35_n_117 | sub_1010_35_n_151));
 assign sub_1010_35_n_166 = ~(n_1352 | ~n_1042);
 assign sub_1010_35_n_165 = ~(sub_1010_35_n_159 | sub_1010_35_n_158);
 assign sub_1010_35_n_164 = ~(sub_1010_35_n_44 & sub_1010_35_n_161);
 assign sub_1010_35_n_163 = ~sub_1010_35_n_162;
 assign sub_1010_35_n_162 = ~(sub_1010_35_n_106 | (sub_1010_35_n_131 | sub_1010_35_n_110));
 assign sub_1010_35_n_157 = ~sub_1010_35_n_44;
 assign sub_1010_35_n_156 = ~(sub_1010_35_n_114 | sub_1010_35_n_138);
 assign sub_1010_35_n_155 = ~(sub_1010_35_n_101 | (sub_1010_35_n_66 & sub_1010_35_n_10));
 assign sub_1010_35_n_161 = ~(sub_1010_35_n_126 | sub_1010_35_n_128);
 assign sub_1010_35_n_160 = ~(sub_1010_35_n_8 & (sub_1010_35_n_6 | sub_1010_35_n_91));
 assign sub_1010_35_n_159 = ~(sub_1010_35_n_141 & sub_1010_35_n_129);
 assign sub_1010_35_n_158 = ~(sub_1010_35_n_119 & sub_1010_35_n_112);
 assign sub_1010_35_n_44 = ~(sub_1010_35_n_18 | sub_1010_35_n_118);
 assign sub_1010_35_n_154 = ~sub_1010_35_n_153;
 assign sub_1010_35_n_152 = ~sub_1010_35_n_151;
 assign sub_1010_35_n_149 = ~sub_1010_35_n_148;
 assign sub_1010_35_n_146 = ~(sub_1010_35_n_77 | (sub_1010_35_n_87 & sub_1010_35_n_74));
 assign sub_1010_35_n_145 = ~(sub_1010_35_n_7 & (sub_1010_35_n_12 | sub_1010_35_n_93));
 assign sub_1010_35_n_144 = ~(sub_1010_35_n_125 | ~sub_1010_35_n_80);
 assign sub_1010_35_n_143 = ~(sub_1010_35_n_4 & (sub_1010_35_n_2 | sub_1010_35_n_58));
 assign sub_1010_35_n_153 = ~(sub_1010_35_n_104 | ~sub_1010_35_n_81);
 assign sub_1010_35_n_151 = ~(sub_1010_35_n_124 | ~sub_1010_35_n_1);
 assign sub_1010_35_n_150 = ~(sub_1010_35_n_14 & (sub_1010_35_n_60 | sub_1010_35_n_75));
 assign sub_1010_35_n_148 = ~(sub_1010_35_n_103 | ~sub_1010_35_n_99);
 assign sub_1010_35_n_147 = ~(sub_1010_35_n_122 | ~sub_1010_35_n_79);
 assign sub_1010_35_n_142 = ~sub_1010_35_n_141;
 assign sub_1010_35_n_139 = ~sub_1010_35_n_20;
 assign sub_1010_35_n_125 = ~(sub_1010_35_n_11 | sub_1010_35_n_86);
 assign sub_1010_35_n_124 = ~(sub_1010_35_n_85 | ~sub_1010_35_n_9);
 assign sub_1010_35_n_123 = ~(sub_1010_35_n_90 | sub_1010_35_n_86);
 assign sub_1010_35_n_122 = ~(sub_1010_35_n_59 | ~sub_1010_35_n_69);
 assign sub_1010_35_n_141 = ~(sub_1010_35_n_96 | sub_1010_35_n_91);
 assign sub_1010_35_n_140 = ~(sub_1010_35_n_2 & sub_1010_35_n_95);
 assign sub_1010_35_n_138 = ~(sub_1010_35_n_3 & sub_1010_35_n_10);
 assign sub_1010_35_n_137 = ~(sub_1010_35_n_60 & sub_1010_35_n_63);
 assign sub_1010_35_n_136 = ~(sub_1010_35_n_98 & sub_1010_35_n_100);
 assign sub_1010_35_n_135 = ~(sub_1010_35_n_6 & sub_1010_35_n_97);
 assign sub_1010_35_n_134 = ~(sub_1010_35_n_43 & sub_1010_35_n_10);
 assign sub_1010_35_n_133 = ~(sub_1010_35_n_37 & sub_1010_35_n_3);
 assign sub_1010_35_n_132 = ~(sub_1010_35_n_99 & sub_1010_35_n_89);
 assign sub_1010_35_n_131 = ~(sub_1010_35_n_100 & ~n_1244);
 assign sub_1010_35_n_130 = ~(sub_1010_35_n_1 & sub_1010_35_n_9);
 assign sub_1010_35_n_129 = ~(sub_1010_35_n_41 | sub_1010_35_n_93);
 assign sub_1010_35_n_128 = ~(sub_1010_35_n_13 & ~sub_1010_35_n_61);
 assign sub_1010_35_n_127 = ~(sub_1010_35_n_85 & sub_1010_35_n_70);
 assign sub_1010_35_n_126 = ~(sub_1010_35_n_92 & ~sub_1010_35_n_65);
 assign sub_1010_35_n_120 = ~sub_1010_35_n_119;
 assign sub_1010_35_n_118 = ~sub_1010_35_n_117;
 assign sub_1010_35_n_111 = ~sub_1010_35_n_110;
 assign sub_1010_35_n_106 = ~sub_1010_35_n_105;
 assign sub_1010_35_n_104 = ~(sub_1010_35_n_64 | sub_1010_35_n_65);
 assign sub_1010_35_n_103 = ~(sub_1010_35_n_40 | sub_1010_35_n_88);
 assign T_5_0_ = ~(sub_1010_35_n_83 & (~{in2[5]} | {in1[0]}));
 assign sub_1010_35_n_121 = ~(sub_1010_35_n_59 & sub_1010_35_n_38);
 assign sub_1010_35_n_119 = ~(sub_1010_35_n_62 | sub_1010_35_n_75);
 assign sub_1010_35_n_117 = ~(sub_1010_35_n_71 | sub_1010_35_n_73);
 assign sub_1010_35_n_116 = ~(sub_1010_35_n_84 & sub_1010_35_n_13);
 assign sub_1010_35_n_115 = ~(sub_1010_35_n_64 & sub_1010_35_n_92);
 assign sub_1010_35_n_114 = ~(sub_1010_35_n_5 & sub_1010_35_n_89);
 assign sub_1010_35_n_113 = ~(sub_1010_35_n_39 & sub_1010_35_n_74);
 assign sub_1010_35_n_112 = ~(sub_1010_35_n_94 | sub_1010_35_n_58);
 assign sub_1010_35_n_110 = ~(sub_1010_35_n_38 & ~sub_1010_35_n_68);
 assign sub_1010_35_n_109 = ~(sub_1010_35_n_42 & sub_1010_35_n_72);
 assign sub_1010_35_n_108 = ~(sub_1010_35_n_78 & sub_1010_35_n_0);
 assign sub_1010_35_n_107 = ~(sub_1010_35_n_79 & sub_1010_35_n_69);
 assign sub_1010_35_n_105 = ~(n_1299 | (n_1363 | (n_832 | n_1275)));
 assign sub_1010_35_n_101 = ~sub_1010_35_n_43;
 assign sub_1010_35_n_100 = ~sub_1010_35_n_82;
 assign sub_1010_35_n_97 = ~sub_1010_35_n_96;
 assign sub_1010_35_n_95 = ~sub_1010_35_n_94;
 assign sub_1010_35_n_89 = ~sub_1010_35_n_88;
 assign sub_1010_35_n_87 = ~sub_1010_35_n_42;
 assign sub_1010_35_n_43 = ~(sub_1010_35_n_50 & R_6_6_);
 assign sub_1010_35_n_82 = ~(R_6_25_ | ~n_1088);
 assign sub_1010_35_n_99 = ~(R_6_4_ & ~n_1051);
 assign sub_1010_35_n_98 = ~(R_6_25_ & ~n_1088);
 assign sub_1010_35_n_96 = ~(R_6_7_ | ~n_1219);
 assign sub_1010_35_n_94 = ~(R_6_13_ | ~n_1184);
 assign sub_1010_35_n_93 = ~(R_6_10_ | ~n_1067);
 assign sub_1010_35_n_92 = ~(sub_1010_35_n_52 & ~sub_1010_35_n_51);
 assign sub_1010_35_n_91 = ~(R_6_8_ | ~n_1164);
 assign sub_1010_35_n_90 = ~(R_6_1_ | ~n_1103);
 assign sub_1010_35_n_88 = ~(R_6_4_ | ~n_1051);
 assign sub_1010_35_n_42 = ~(R_6_17_ & ~n_1033);
 assign sub_1010_35_n_41 = ~(R_6_9_ | ~n_1347);
 assign sub_1010_35_n_40 = ~(sub_1010_35_n_57 & R_6_3_);
 assign sub_1010_35_n_86 = ~(R_6_2_ | ~n_1115);
 assign sub_1010_35_n_85 = ~(R_6_15_ & ~n_1138);
 assign sub_1010_35_n_84 = ~(R_6_21_ & ~n_1179);
 assign sub_1010_35_n_83 = ~({in1[0]} & ~{in2[5]});
 assign sub_1010_35_n_77 = ~sub_1010_35_n_39;
 assign sub_1010_35_n_74 = ~sub_1010_35_n_73;
 assign sub_1010_35_n_72 = ~sub_1010_35_n_71;
 assign sub_1010_35_n_69 = ~sub_1010_35_n_68;
 assign sub_1010_35_n_38 = ~sub_1010_35_n_67;
 assign sub_1010_35_n_66 = ~sub_1010_35_n_37;
 assign sub_1010_35_n_63 = ~sub_1010_35_n_62;
 assign sub_1010_35_n_81 = ~(R_6_20_ & ~n_1368);
 assign sub_1010_35_n_80 = ~(R_6_2_ & ~n_1115);
 assign sub_1010_35_n_79 = ~(R_6_24_ & ~n_1373);
 assign sub_1010_35_n_78 = ~(sub_1010_35_n_54 & R_6_0_);
 assign sub_1010_35_n_39 = ~(R_6_18_ & ~n_1304);
 assign sub_1010_35_n_76 = ~(R_6_22_ & ~n_1294);
 assign sub_1010_35_n_75 = ~(R_6_12_ | ~n_1261);
 assign sub_1010_35_n_73 = ~(R_6_18_ | ~n_1304);
 assign sub_1010_35_n_71 = ~(R_6_17_ | ~n_1033);
 assign sub_1010_35_n_70 = ~(sub_1010_35_n_53 & ~sub_1010_35_n_55);
 assign sub_1010_35_n_68 = ~(R_6_24_ | ~n_1373);
 assign sub_1010_35_n_67 = ~(R_6_23_ | ~n_1061);
 assign sub_1010_35_n_37 = ~(sub_1010_35_n_56 & R_6_5_);
 assign sub_1010_35_n_65 = ~(R_6_20_ | ~n_1368);
 assign sub_1010_35_n_64 = ~(sub_1010_35_n_51 & R_6_19_);
 assign sub_1010_35_n_62 = ~(R_6_11_ | ~n_1028);
 assign sub_1010_35_n_61 = ~(R_6_22_ | ~n_1294);
 assign sub_1010_35_n_60 = ~(R_6_11_ & ~n_1028);
 assign sub_1010_35_n_59 = ~(R_6_23_ & ~n_1061);
 assign sub_1010_35_n_58 = ~(R_6_14_ | ~n_1093);
 assign sub_1010_35_n_57 = ~n_1342;
 assign sub_1010_35_n_56 = ~n_1098;
 assign sub_1010_35_n_55 = ~n_1138;
 assign sub_1010_35_n_54 = ~n_1352;
 assign sub_1010_35_n_53 = ~R_6_15_;
 assign sub_1010_35_n_52 = ~R_6_19_;
 assign sub_1010_35_n_51 = ~n_1214;
 assign sub_1010_35_n_50 = ~n_1169;
 assign sub_1010_35_n_49 = ~R_6_16_;
 assign sub_1010_35_n_36 = (sub_1010_35_n_76 & (sub_1010_35_n_84 | sub_1010_35_n_61));
 assign sub_1010_35_n_35 = ~(sub_1010_35_n_2 & ~(sub_1010_35_n_95 & sub_1010_35_n_221));
 assign sub_1010_35_n_34 = ~(sub_1010_35_n_60 & ~(sub_1010_35_n_63 & sub_1010_35_n_33));
 assign sub_1010_35_n_33 = ~(sub_1010_35_n_195 & sub_1010_35_n_169);
 assign sub_1010_35_n_32 = ~(sub_1010_35_n_151 & (sub_1010_35_n_18 | sub_1010_35_n_202));
 assign sub_1010_35_n_31 = ~(sub_1010_35_n_157 | sub_1010_35_n_126);
 assign sub_1010_35_n_30 = ~(sub_1010_35_n_148 & (sub_1010_35_n_114 | sub_1010_35_n_186));
 assign sub_1010_35_n_29 = (sub_1010_35_n_98 | n_1244);
 assign sub_1010_35_n_28 = ~(sub_1010_35_n_7 & ~sub_1010_35_n_93);
 assign sub_1010_35_n_27 = ~(sub_1010_35_n_8 & ~sub_1010_35_n_91);
 assign sub_1010_35_n_26 = ~(sub_1010_35_n_11 & ~sub_1010_35_n_90);
 assign sub_1010_35_n_25 = ~(sub_1010_35_n_12 & (sub_1010_35_n_41 | sub_1010_35_n_205));
 assign sub_1010_35_n_24 = ~(sub_1010_35_n_184 & sub_1010_35_n_11);
 assign sub_1010_35_n_23 = (sub_1010_35_n_40 & sub_1010_35_n_5);
 assign sub_1010_35_n_22 = ~(sub_1010_35_n_80 & ~sub_1010_35_n_86);
 assign sub_1010_35_n_21 = ~(sub_1010_35_n_84 & (~sub_1010_35_n_13 | sub_1010_35_n_206));
 assign sub_1010_35_n_20 = ~(sub_1010_35_n_14 & ~sub_1010_35_n_75);
 assign sub_1010_35_n_19 = ~(sub_1010_35_n_41 | ~sub_1010_35_n_12);
 assign sub_1010_35_n_18 = ~(sub_1010_35_n_70 & sub_1010_35_n_9);
 assign sub_1010_35_n_17 = ~(sub_1010_35_n_81 & ~sub_1010_35_n_65);
 assign sub_1010_35_n_16 = ~(sub_1010_35_n_76 & ~sub_1010_35_n_61);
 assign sub_1010_35_n_15 = ~(sub_1010_35_n_4 & ~sub_1010_35_n_58);
 assign sub_1010_35_n_14 = ~(R_6_12_ & ~n_1261);
 assign sub_1010_35_n_13 = ~(n_1179 & ~R_6_21_);
 assign sub_1010_35_n_12 = ~(R_6_9_ & ~n_1347);
 assign sub_1010_35_n_11 = ~(R_6_1_ & ~n_1103);
 assign sub_1010_35_n_10 = (R_6_6_ | sub_1010_35_n_50);
 assign sub_1010_35_n_9 = ~(sub_1010_35_n_49 & n_1174);
 assign sub_1010_35_n_8 = ~(R_6_8_ & ~n_1164);
 assign sub_1010_35_n_7 = ~(R_6_10_ & ~n_1067);
 assign sub_1010_35_n_6 = ~(R_6_7_ & ~n_1219);
 assign sub_1010_35_n_5 = (R_6_3_ | sub_1010_35_n_57);
 assign sub_1010_35_n_4 = ~(R_6_14_ & ~n_1093);
 assign sub_1010_35_n_3 = (R_6_5_ | sub_1010_35_n_56);
 assign sub_1010_35_n_2 = ~(R_6_13_ & ~n_1184);
 assign sub_1010_35_n_1 = (sub_1010_35_n_49 | n_1174);
 assign sub_1010_35_n_0 = (R_6_0_ | sub_1010_35_n_54);
 assign T_4_27_ = ((sub_1040_34_n_21 & sub_1040_34_n_29) | ~(sub_1040_34_n_21 | sub_1040_34_n_29));
 assign T_4_15_ = ((sub_1040_34_n_139 & ~sub_1040_34_n_33) | (sub_1040_34_n_26 & sub_1040_34_n_33));
 assign T_4_26_ = ((sub_1040_34_n_228 & sub_1040_34_n_28) | ~(sub_1040_34_n_228 | sub_1040_34_n_28));
 assign T_4_25_ = ((sub_1040_34_n_232 & sub_1040_34_n_22) | ~(sub_1040_34_n_232 | sub_1040_34_n_22));
 assign T_4_23_ = ((sub_1040_34_n_231 & sub_1040_34_n_32) | ~(sub_1040_34_n_231 | sub_1040_34_n_32));
 assign T_4_21_ = ((sub_1040_34_n_230 & n_876) | ~(sub_1040_34_n_230 | n_876));
 assign T_4_19_ = ((sub_1040_34_n_229 & sub_1040_34_n_30) | ~(sub_1040_34_n_229 | sub_1040_34_n_30));
 assign T_4_18_ = ((sub_1040_34_n_50 & sub_1040_34_n_132) | ~(sub_1040_34_n_50 | sub_1040_34_n_132));
 assign sub_1040_34_n_232 = ~(sub_1040_34_n_78 | (~sub_1040_34_n_73 & sub_1040_34_n_214));
 assign sub_1040_34_n_231 = ~(n_859 & (~sub_1040_34_n_3 | sub_1040_34_n_215));
 assign sub_1040_34_n_230 = ~(sub_1040_34_n_72 | (~sub_1040_34_n_100 & sub_1040_34_n_212));
 assign sub_1040_34_n_229 = ~(n_852 | (~n_848 & sub_1040_34_n_39));
 assign sub_1040_34_n_228 = ~(sub_1040_34_n_147 | (~sub_1040_34_n_137 & sub_1040_34_n_214));
 assign T_4_20_ = ((sub_1040_34_n_212 & sub_1040_34_n_121) | ~(sub_1040_34_n_212 | sub_1040_34_n_121));
 assign T_4_14_ = ~((sub_1040_34_n_216 | sub_1040_34_n_20) & ~(sub_1040_34_n_216 & sub_1040_34_n_20));
 assign T_4_13_ = ~((sub_1040_34_n_219 | sub_1040_34_n_24) & ~(sub_1040_34_n_219 & sub_1040_34_n_24));
 assign T_4_11_ = ~((sub_1040_34_n_217 | sub_1040_34_n_35) & ~(sub_1040_34_n_217 & sub_1040_34_n_35));
 assign T_4_24_ = ((sub_1040_34_n_214 & sub_1040_34_n_127) | ~(sub_1040_34_n_214 | sub_1040_34_n_127));
 assign T_4_22_ = ((sub_1040_34_n_215 & sub_1040_34_n_34) | ~(sub_1040_34_n_215 | sub_1040_34_n_34));
 assign T_4_17_ = ((sub_1040_34_n_218 & sub_1040_34_n_141) | ~(sub_1040_34_n_218 | sub_1040_34_n_141));
 assign T_4_32_ = ~(sub_1040_34_n_204 | sub_1040_34_n_185);
 assign sub_1040_34_n_219 = ~(sub_1040_34_n_76 | (~n_893 & sub_1040_34_n_41));
 assign sub_1040_34_n_218 = ~(n_860 | (~sub_1040_34_n_85 & sub_1040_34_n_199));
 assign sub_1040_34_n_217 = ~(sub_1040_34_n_94 | (~n_840 & sub_1040_34_n_202));
 assign sub_1040_34_n_216 = ~(sub_1040_34_n_150 | (~sub_1040_34_n_125 & sub_1040_34_n_41));
 assign sub_1040_34_n_215 = ~(sub_1040_34_n_42 | (~sub_1040_34_n_163 & sub_1040_34_n_199));
 assign sub_1040_34_n_214 = ~(sub_1040_34_n_205 & ~sub_1040_34_n_179);
 assign sub_1040_34_n_50 = ~sub_1040_34_n_39;
 assign T_4_16_ = ~((sub_1040_34_n_200 | sub_1040_34_n_140) & ~(sub_1040_34_n_200 & sub_1040_34_n_140));
 assign T_4_7_ = ((sub_1040_34_n_197 & sub_1040_34_n_36) | ~(sub_1040_34_n_197 | sub_1040_34_n_36));
 assign T_4_12_ = ((sub_1040_34_n_41 & sub_1040_34_n_19) | ~(sub_1040_34_n_41 | sub_1040_34_n_19));
 assign T_4_10_ = ~((sub_1040_34_n_203 | sub_1040_34_n_118) & ~(sub_1040_34_n_203 & sub_1040_34_n_118));
 assign T_4_9_ = ((sub_1040_34_n_201 & sub_1040_34_n_37) | ~(sub_1040_34_n_201 | sub_1040_34_n_37));
 assign sub_1040_34_n_212 = ~(sub_1040_34_n_40 & ~sub_1040_34_n_171);
 assign sub_1040_34_n_206 = ~(sub_1040_34_n_199 & ~sub_1040_34_n_133);
 assign sub_1040_34_n_205 = ~(sub_1040_34_n_199 & ~sub_1040_34_n_164);
 assign sub_1040_34_n_204 = ~(sub_1040_34_n_198 | ~sub_1040_34_n_173);
 assign sub_1040_34_n_203 = ~sub_1040_34_n_202;
 assign sub_1040_34_n_202 = ~(sub_1040_34_n_193 & ~sub_1040_34_n_160);
 assign sub_1040_34_n_201 = ~(sub_1040_34_n_103 | (~n_874 & sub_1040_34_n_190));
 assign sub_1040_34_n_200 = ~sub_1040_34_n_199;
 assign sub_1040_34_n_199 = ~sub_1040_34_n_198;
 assign sub_1040_34_n_198 = ~(sub_1040_34_n_192 | sub_1040_34_n_177);
 assign sub_1040_34_n_197 = ~(sub_1040_34_n_67 & (~n_885 | sub_1040_34_n_191));
 assign T_4_5_ = ~((sub_1040_34_n_188 | sub_1040_34_n_126) & ~(sub_1040_34_n_188 & sub_1040_34_n_126));
 assign T_4_8_ = ~((sub_1040_34_n_190 | sub_1040_34_n_27) & ~(sub_1040_34_n_190 & sub_1040_34_n_27));
 assign sub_1040_34_n_194 = ~(sub_1040_34_n_190 & ~sub_1040_34_n_157);
 assign sub_1040_34_n_193 = ~(sub_1040_34_n_190 & ~sub_1040_34_n_123);
 assign sub_1040_34_n_192 = ~(sub_1040_34_n_189 | ~sub_1040_34_n_162);
 assign sub_1040_34_n_191 = ~(sub_1040_34_n_149 | (~sub_1040_34_n_138 & n_897));
 assign sub_1040_34_n_190 = ~sub_1040_34_n_189;
 assign sub_1040_34_n_189 = ~(sub_1040_34_n_170 | (n_897 & sub_1040_34_n_154));
 assign sub_1040_34_n_188 = ~(sub_1040_34_n_87 & (~n_899 | sub_1040_34_n_184));
 assign T_4_4_ = ((sub_1040_34_n_184 & sub_1040_34_n_25) | ~(sub_1040_34_n_184 | sub_1040_34_n_25));
 assign T_4_3_ = ((sub_1040_34_n_182 & sub_1040_34_n_128) | ~(sub_1040_34_n_182 | sub_1040_34_n_128));
 assign sub_1040_34_n_185 = ~(sub_1040_34_n_175 & (sub_1040_34_n_178 | sub_1040_34_n_161));
 assign sub_1040_34_n_184 = ~n_897;
 assign sub_1040_34_n_183 = ~(sub_1040_34_n_176 & sub_1040_34_n_145);
 assign sub_1040_34_n_182 = ~(sub_1040_34_n_180 & ~sub_1040_34_n_13);
 assign T_4_2_ = ~((sub_1040_34_n_174 | sub_1040_34_n_31) & ~(sub_1040_34_n_174 & sub_1040_34_n_31));
 assign sub_1040_34_n_180 = ~(sub_1040_34_n_174 & ~sub_1040_34_n_104);
 assign sub_1040_34_n_179 = ~sub_1040_34_n_178;
 assign sub_1040_34_n_178 = ~(sub_1040_34_n_169 | (sub_1040_34_n_171 & sub_1040_34_n_158));
 assign sub_1040_34_n_177 = ~(sub_1040_34_n_168 & (sub_1040_34_n_167 | sub_1040_34_n_159));
 assign sub_1040_34_n_176 = ~(sub_1040_34_n_174 & sub_1040_34_n_130);
 assign sub_1040_34_n_175 = ~(n_834 & (sub_1040_34_n_146 | (sub_1040_34_n_147 & sub_1040_34_n_134)));
 assign sub_1040_34_n_174 = ~(sub_1040_34_n_165 & (sub_1040_34_n_166 & sub_1040_34_n_111));
 assign sub_1040_34_n_173 = ~(sub_1040_34_n_161 | sub_1040_34_n_164);
 assign T_4_1_ = ((sub_1040_34_n_119 & n_1132) | ~(sub_1040_34_n_119 | n_1132));
 assign sub_1040_34_n_171 = ~(sub_1040_34_n_153 & (~sub_1040_34_n_136 | sub_1040_34_n_152));
 assign sub_1040_34_n_170 = ~(sub_1040_34_n_156 & (sub_1040_34_n_148 | sub_1040_34_n_131));
 assign sub_1040_34_n_169 = ~(sub_1040_34_n_45 & (n_904 | sub_1040_34_n_120));
 assign sub_1040_34_n_168 = ~(sub_1040_34_n_144 | (sub_1040_34_n_150 & sub_1040_34_n_129));
 assign sub_1040_34_n_167 = ~(sub_1040_34_n_143 | (sub_1040_34_n_160 & sub_1040_34_n_142));
 assign sub_1040_34_n_166 = ~(n_1132 & R_5_0_);
 assign sub_1040_34_n_165 = ~(n_1132 & ~n_1352);
 assign sub_1040_34_n_164 = ~(sub_1040_34_n_38 & sub_1040_34_n_158);
 assign sub_1040_34_n_163 = ~(sub_1040_34_n_38 & sub_1040_34_n_115);
 assign sub_1040_34_n_162 = ~(sub_1040_34_n_157 | sub_1040_34_n_159);
 assign sub_1040_34_n_161 = ~(sub_1040_34_n_155 & sub_1040_34_n_134);
 assign sub_1040_34_n_156 = ~(n_881 | (n_887 & n_882));
 assign sub_1040_34_n_155 = ~(sub_1040_34_n_117 | sub_1040_34_n_137);
 assign sub_1040_34_n_154 = ~(sub_1040_34_n_138 | sub_1040_34_n_131);
 assign sub_1040_34_n_153 = ~(n_844 | (n_852 & sub_1040_34_n_102));
 assign sub_1040_34_n_160 = ~(n_905 & (n_877 | n_866));
 assign sub_1040_34_n_159 = ~(sub_1040_34_n_124 & sub_1040_34_n_129);
 assign sub_1040_34_n_158 = ~(sub_1040_34_n_114 | sub_1040_34_n_120);
 assign sub_1040_34_n_157 = ~(sub_1040_34_n_122 & sub_1040_34_n_142);
 assign sub_1040_34_n_149 = ~sub_1040_34_n_148;
 assign sub_1040_34_n_146 = ~(sub_1040_34_n_90 & (sub_1040_34_n_4 | sub_1040_34_n_99));
 assign sub_1040_34_n_145 = ~(sub_1040_34_n_88 | (sub_1040_34_n_13 & sub_1040_34_n_80));
 assign sub_1040_34_n_144 = ~(sub_1040_34_n_14 & (n_878 | n_845));
 assign sub_1040_34_n_143 = ~(n_906 & (n_839 | n_892));
 assign sub_1040_34_n_152 = ~(n_851 | (~n_850 & n_860));
 assign sub_1040_34_n_151 = ~(sub_1040_34_n_113 | ~sub_1040_34_n_91);
 assign sub_1040_34_n_150 = ~(n_863 & (n_891 | n_865));
 assign sub_1040_34_n_148 = ~(sub_1040_34_n_92 | (n_900 & n_884));
 assign sub_1040_34_n_147 = ~(sub_1040_34_n_89 & (sub_1040_34_n_77 | sub_1040_34_n_86));
 assign sub_1040_34_n_139 = ~sub_1040_34_n_26;
 assign sub_1040_34_n_130 = ~(sub_1040_34_n_104 | sub_1040_34_n_79);
 assign sub_1040_34_n_142 = ~(n_840 | n_892);
 assign sub_1040_34_n_141 = ~(n_851 | n_850);
 assign sub_1040_34_n_140 = ~(n_860 | sub_1040_34_n_85);
 assign sub_1040_34_n_138 = ~(n_899 & n_884);
 assign sub_1040_34_n_137 = ~(sub_1040_34_n_74 & ~n_858);
 assign sub_1040_34_n_136 = ~(n_848 | n_847);
 assign sub_1040_34_n_135 = ~(sub_1040_34_n_67 & n_885);
 assign sub_1040_34_n_134 = ~(sub_1040_34_n_82 | sub_1040_34_n_99);
 assign sub_1040_34_n_133 = ~(sub_1040_34_n_15 & ~n_850);
 assign sub_1040_34_n_132 = ~(n_852 | n_848);
 assign sub_1040_34_n_131 = ~(n_885 & n_882);
 assign sub_1040_34_n_125 = ~sub_1040_34_n_124;
 assign sub_1040_34_n_123 = ~sub_1040_34_n_122;
 assign sub_1040_34_n_117 = ~n_834;
 assign sub_1040_34_n_115 = ~sub_1040_34_n_114;
 assign sub_1040_34_n_113 = ~(sub_1040_34_n_71 | ~sub_1040_34_n_64);
 assign T_4_0_ = ~(sub_1040_34_n_93 & (~{in2[4]} | {in1[0]}));
 assign sub_1040_34_n_129 = ~(n_864 | n_845);
 assign sub_1040_34_n_128 = ~(sub_1040_34_n_1 & sub_1040_34_n_80);
 assign sub_1040_34_n_127 = ~(sub_1040_34_n_77 & sub_1040_34_n_74);
 assign sub_1040_34_n_126 = ~(n_886 & n_884);
 assign sub_1040_34_n_124 = ~(n_893 | n_865);
 assign sub_1040_34_n_122 = ~(n_874 | n_866);
 assign sub_1040_34_n_121 = ~(n_857 & sub_1040_34_n_5);
 assign sub_1040_34_n_120 = ~(sub_1040_34_n_3 & ~n_868);
 assign sub_1040_34_n_119 = ~(sub_1040_34_n_111 & sub_1040_34_n_0);
 assign sub_1040_34_n_118 = ~(sub_1040_34_n_94 | n_840);
 assign sub_1040_34_n_116 = ~(n_1299 | (n_1363 | (n_832 | n_1275)));
 assign sub_1040_34_n_114 = ~(sub_1040_34_n_5 & ~n_896);
 assign sub_1040_34_n_49 = ~sub_1040_34_n_108;
 assign sub_1040_34_n_103 = ~n_877;
 assign sub_1040_34_n_102 = ~n_847;
 assign sub_1040_34_n_100 = ~sub_1040_34_n_5;
 assign sub_1040_34_n_94 = ~n_839;
 assign sub_1040_34_n_111 = ~(sub_1040_34_n_60 & R_5_0_);
 assign sub_1040_34_n_110 = ~(n_1169 | sub_1040_34_n_54);
 assign sub_1040_34_n_109 = ~(R_5_22_ & ~n_1294);
 assign sub_1040_34_n_108 = ~(R_5_15_ & ~n_1138);
 assign sub_1040_34_n_107 = ~(sub_1040_34_n_61 & ~sub_1040_34_n_59);
 assign sub_1040_34_n_106 = ~(R_5_13_ | ~n_1184);
 assign sub_1040_34_n_105 = ~(R_5_22_ | ~n_1294);
 assign sub_1040_34_n_104 = ~(R_5_1_ | ~n_1103);
 assign sub_1040_34_n_48 = ~(R_5_7_ & ~n_1219);
 assign sub_1040_34_n_101 = ~(R_5_18_ | ~n_1304);
 assign sub_1040_34_n_99 = ~(n_870 | ~n_1245);
 assign sub_1040_34_n_98 = ~(R_5_7_ | ~n_1219);
 assign sub_1040_34_n_97 = ~(R_5_14_ | ~n_1093);
 assign sub_1040_34_n_96 = ~(R_5_10_ | ~n_1067);
 assign sub_1040_34_n_95 = ~(R_5_12_ | ~n_1261);
 assign sub_1040_34_n_47 = ~(R_5_21_ & ~n_1179);
 assign sub_1040_34_n_93 = ~({in1[0]} & ~{in2[4]});
 assign sub_1040_34_n_92 = ~n_886;
 assign sub_1040_34_n_88 = ~sub_1040_34_n_1;
 assign sub_1040_34_n_87 = ~n_900;
 assign sub_1040_34_n_85 = ~sub_1040_34_n_15;
 assign sub_1040_34_n_80 = ~sub_1040_34_n_79;
 assign sub_1040_34_n_78 = ~sub_1040_34_n_77;
 assign sub_1040_34_n_76 = ~n_891;
 assign sub_1040_34_n_73 = ~sub_1040_34_n_74;
 assign sub_1040_34_n_72 = ~n_857;
 assign sub_1040_34_n_67 = ~n_887;
 assign sub_1040_34_n_46 = ~(sub_1040_34_n_59 & R_5_4_);
 assign sub_1040_34_n_91 = ~(R_5_20_ & ~n_1368);
 assign sub_1040_34_n_90 = ~(n_870 & ~n_1245);
 assign sub_1040_34_n_89 = ~(sub_1040_34_n_52 & n_855);
 assign sub_1040_34_n_65 = ~(R_5_24_ | ~n_1373);
 assign sub_1040_34_n_86 = ~(n_855 | ~n_1374);
 assign sub_1040_34_n_84 = ~(R_5_9_ | ~n_1347);
 assign sub_1040_34_n_83 = ~(R_5_8_ | ~n_1164);
 assign sub_1040_34_n_82 = ~(n_875 | ~n_1089);
 assign sub_1040_34_n_81 = ~(R_5_17_ | ~n_1033);
 assign sub_1040_34_n_79 = ~(R_5_2_ | ~n_1115);
 assign sub_1040_34_n_77 = ~(sub_1040_34_n_57 & ~n_1062);
 assign sub_1040_34_n_64 = ~(sub_1040_34_n_53 & ~sub_1040_34_n_58);
 assign sub_1040_34_n_75 = ~(R_5_20_ | ~n_1368);
 assign sub_1040_34_n_74 = ~(sub_1040_34_n_56 & ~n_1063);
 assign sub_1040_34_n_71 = ~(R_5_19_ & ~n_1214);
 assign sub_1040_34_n_70 = ~(R_5_11_ | ~n_1028);
 assign sub_1040_34_n_69 = ~(R_5_16_ | ~n_1174);
 assign sub_1040_34_n_68 = ~(n_1033 | sub_1040_34_n_63);
 assign sub_1040_34_n_66 = ~(n_1098 | sub_1040_34_n_55);
 assign sub_1040_34_n_63 = ~R_5_17_;
 assign sub_1040_34_n_62 = ~n_1061;
 assign sub_1040_34_n_61 = ~R_5_4_;
 assign sub_1040_34_n_60 = ~n_1352;
 assign sub_1040_34_n_59 = ~n_1051;
 assign sub_1040_34_n_58 = ~n_1368;
 assign sub_1040_34_n_57 = ~sub_1040_34_n_56;
 assign sub_1040_34_n_56 = ~n_871;
 assign sub_1040_34_n_55 = ~R_5_5_;
 assign sub_1040_34_n_54 = ~R_5_6_;
 assign sub_1040_34_n_53 = ~R_5_20_;
 assign sub_1040_34_n_52 = ~n_1374;
 assign sub_1040_34_n_45 = (n_869 & (n_859 | n_868));
 assign sub_1040_34_n_44 = ~(n_1304 | ~R_5_18_);
 assign T_4_6_ = (sub_1040_34_n_191 ^ sub_1040_34_n_135);
 assign sub_1040_34_n_42 = ~(n_904 & ~(sub_1040_34_n_115 & sub_1040_34_n_171));
 assign sub_1040_34_n_41 = ~(sub_1040_34_n_194 & sub_1040_34_n_167);
 assign sub_1040_34_n_40 = ~(sub_1040_34_n_199 & sub_1040_34_n_38);
 assign sub_1040_34_n_39 = ~(sub_1040_34_n_206 & sub_1040_34_n_152);
 assign sub_1040_34_n_38 = ~(sub_1040_34_n_133 | ~sub_1040_34_n_136);
 assign sub_1040_34_n_37 = ~(n_866 | ~n_905);
 assign sub_1040_34_n_36 = ~(n_882 & ~n_881);
 assign sub_1040_34_n_35 = ~(n_892 | ~n_906);
 assign sub_1040_34_n_34 = (n_859 & sub_1040_34_n_3);
 assign sub_1040_34_n_33 = ~(n_878 & (n_864 | sub_1040_34_n_216));
 assign sub_1040_34_n_32 = ~(n_869 & ~n_868);
 assign sub_1040_34_n_31 = (sub_1040_34_n_13 | sub_1040_34_n_104);
 assign sub_1040_34_n_30 = ~(n_844 | ~sub_1040_34_n_102);
 assign sub_1040_34_n_29 = ~(sub_1040_34_n_90 & ~sub_1040_34_n_99);
 assign sub_1040_34_n_28 = ~(sub_1040_34_n_82 | ~sub_1040_34_n_4);
 assign sub_1040_34_n_27 = ~(n_877 & ~n_874);
 assign sub_1040_34_n_26 = ~(sub_1040_34_n_14 & ~n_845);
 assign sub_1040_34_n_25 = ~(n_900 | ~n_899);
 assign sub_1040_34_n_24 = ~(n_865 | ~n_863);
 assign sub_1040_34_n_23 = ~(sub_1040_34_n_75 | ~sub_1040_34_n_91);
 assign sub_1040_34_n_22 = ~(sub_1040_34_n_86 | ~sub_1040_34_n_89);
 assign sub_1040_34_n_21 = ~(sub_1040_34_n_4 & (sub_1040_34_n_82 | sub_1040_34_n_228));
 assign sub_1040_34_n_20 = ~(n_864 | ~n_878);
 assign sub_1040_34_n_19 = ~(n_891 & ~n_893);
 assign sub_1040_34_n_18 = ~(R_5_10_ & ~n_1067);
 assign sub_1040_34_n_17 = ~(R_5_13_ & ~n_1184);
 assign sub_1040_34_n_16 = ~(R_5_8_ & ~n_1164);
 assign sub_1040_34_n_15 = ~(n_1139 & ~n_853);
 assign sub_1040_34_n_14 = ~(n_842 & ~n_1094);
 assign sub_1040_34_n_13 = ~(n_1103 | ~R_5_1_);
 assign sub_1040_34_n_12 = ~(sub_1040_34_n_55 & n_1098);
 assign sub_1040_34_n_11 = ~(n_1342 & ~R_5_3_);
 assign sub_1040_34_n_10 = ~(n_1342 | ~R_5_3_);
 assign sub_1040_34_n_9 = ~(n_1174 | ~R_5_16_);
 assign sub_1040_34_n_8 = ~(sub_1040_34_n_54 & n_1169);
 assign sub_1040_34_n_7 = ~(R_5_11_ & ~n_1028);
 assign sub_1040_34_n_6 = ~(R_5_9_ & ~n_1347);
 assign sub_1040_34_n_5 = ~(n_1215 & ~n_854);
 assign sub_1040_34_n_4 = ~(n_875 & ~n_1089);
 assign sub_1040_34_n_3 = ~(n_1180 & ~n_856);
 assign sub_1040_34_n_2 = ~(R_5_12_ & ~n_1261);
 assign sub_1040_34_n_1 = ~(R_5_2_ & ~n_1115);
 assign sub_1040_34_n_0 = (R_5_0_ | sub_1040_34_n_60);
 assign T_3_28_ = ~((sub_1070_33_n_238 | sub_1070_33_n_28) & ~(sub_1070_33_n_238 & sub_1070_33_n_28));
 assign T_3_19_ = ~((sub_1070_33_n_236 | sub_1070_33_n_139) & ~(sub_1070_33_n_236 & sub_1070_33_n_139));
 assign T_3_27_ = ((sub_1070_33_n_23 & sub_1070_33_n_33) | ~(sub_1070_33_n_23 | sub_1070_33_n_33));
 assign T_3_25_ = ~((sub_1070_33_n_237 | sub_1070_33_n_29) & ~(sub_1070_33_n_237 & sub_1070_33_n_29));
 assign T_3_23_ = ((sub_1070_33_n_24 & sub_1070_33_n_34) | ~(sub_1070_33_n_24 | sub_1070_33_n_34));
 assign T_3_21_ = ((sub_1070_33_n_49 & sub_1070_33_n_142) | ~(sub_1070_33_n_49 | sub_1070_33_n_142));
 assign T_3_18_ = ~((sub_1070_33_n_224 | sub_1070_33_n_25) & ~(sub_1070_33_n_224 & sub_1070_33_n_25));
 assign sub_1070_33_n_238 = ~(sub_1070_33_n_178 | (sub_1070_33_n_223 & sub_1070_33_n_164));
 assign sub_1070_33_n_237 = ~(sub_1070_33_n_102 | (sub_1070_33_n_223 & sub_1070_33_n_99));
 assign sub_1070_33_n_236 = ~(sub_1070_33_n_77 | (~sub_1070_33_n_78 & sub_1070_33_n_224));
 assign T_3_22_ = ~((sub_1070_33_n_48 | sub_1070_33_n_35) & ~(sub_1070_33_n_48 & sub_1070_33_n_35));
 assign T_3_14_ = ~((sub_1070_33_n_41 | sub_1070_33_n_111) & ~(sub_1070_33_n_41 & sub_1070_33_n_111));
 assign T_3_13_ = ((sub_1070_33_n_225 & sub_1070_33_n_131) | ~(sub_1070_33_n_225 | sub_1070_33_n_131));
 assign T_3_11_ = ~((sub_1070_33_n_39 | sub_1070_33_n_128) & ~(sub_1070_33_n_39 & sub_1070_33_n_128));
 assign T_3_26_ = ((sub_1070_33_n_220 & sub_1070_33_n_31) | ~(sub_1070_33_n_220 | sub_1070_33_n_31));
 assign T_3_24_ = ~((sub_1070_33_n_223 | sub_1070_33_n_116) & ~(sub_1070_33_n_223 & sub_1070_33_n_116));
 assign T_3_17_ = ((sub_1070_33_n_132 & ~sub_1070_33_n_221) | (sub_1070_33_n_133 & sub_1070_33_n_221));
 assign T_3_20_ = ((sub_1070_33_n_214 & sub_1070_33_n_141) | ~(sub_1070_33_n_214 | sub_1070_33_n_141));
 assign T_3_32_ = ~sub_1070_33_n_222;
 assign sub_1070_33_n_222 = ~(sub_1070_33_n_212 & sub_1070_33_n_199);
 assign sub_1070_33_n_225 = ~(sub_1070_33_n_70 | (~sub_1070_33_n_71 & sub_1070_33_n_210));
 assign sub_1070_33_n_221 = ~(sub_1070_33_n_108 | (~sub_1070_33_n_81 & sub_1070_33_n_206));
 assign sub_1070_33_n_224 = ~(sub_1070_33_n_42 & ~sub_1070_33_n_166);
 assign sub_1070_33_n_223 = ~(sub_1070_33_n_213 & ~sub_1070_33_n_190);
 assign T_3_9_ = ~((sub_1070_33_n_208 | sub_1070_33_n_121) & ~(sub_1070_33_n_208 & sub_1070_33_n_121));
 assign T_3_10_ = ~((sub_1070_33_n_209 | sub_1070_33_n_117) & ~(sub_1070_33_n_209 & sub_1070_33_n_117));
 assign T_3_12_ = ((sub_1070_33_n_211 & sub_1070_33_n_129) | ~(sub_1070_33_n_211 | sub_1070_33_n_129));
 assign T_3_7_ = ((sub_1070_33_n_207 & sub_1070_33_n_140) | ~(sub_1070_33_n_207 | sub_1070_33_n_140));
 assign T_3_16_ = ~((sub_1070_33_n_206 | sub_1070_33_n_27) & ~(sub_1070_33_n_206 & sub_1070_33_n_27));
 assign sub_1070_33_n_220 = ~(sub_1070_33_n_47 | (sub_1070_33_n_206 & sub_1070_33_n_180));
 assign sub_1070_33_n_214 = ~(sub_1070_33_n_202 & ~sub_1070_33_n_183);
 assign sub_1070_33_n_213 = ~(sub_1070_33_n_206 & ~sub_1070_33_n_168);
 assign sub_1070_33_n_212 = ~(sub_1070_33_n_206 & ~sub_1070_33_n_181);
 assign sub_1070_33_n_210 = ~sub_1070_33_n_211;
 assign sub_1070_33_n_211 = ~(sub_1070_33_n_45 | (~sub_1070_33_n_160 & sub_1070_33_n_197));
 assign sub_1070_33_n_209 = ~sub_1070_33_n_46;
 assign sub_1070_33_n_208 = ~(sub_1070_33_n_5 | (~sub_1070_33_n_72 & sub_1070_33_n_196));
 assign sub_1070_33_n_207 = ~(sub_1070_33_n_87 | (~sub_1070_33_n_67 & sub_1070_33_n_198));
 assign sub_1070_33_n_206 = ~(sub_1070_33_n_201 & sub_1070_33_n_185);
 assign T_3_6_ = ((sub_1070_33_n_198 & sub_1070_33_n_22) | ~(sub_1070_33_n_198 | sub_1070_33_n_22));
 assign T_3_5_ = ~((sub_1070_33_n_26 | sub_1070_33_n_37) & ~(sub_1070_33_n_26 & sub_1070_33_n_37));
 assign T_3_8_ = ((sub_1070_33_n_196 & sub_1070_33_n_36) | ~(sub_1070_33_n_196 | sub_1070_33_n_36));
 assign sub_1070_33_n_202 = ~(sub_1070_33_n_200 | sub_1070_33_n_192);
 assign sub_1070_33_n_201 = ~(sub_1070_33_n_197 & sub_1070_33_n_169);
 assign sub_1070_33_n_200 = ~(sub_1070_33_n_195 | sub_1070_33_n_179);
 assign sub_1070_33_n_199 = ~(sub_1070_33_n_184 | (sub_1070_33_n_190 & sub_1070_33_n_170));
 assign sub_1070_33_n_198 = ~(sub_1070_33_n_153 & (~sub_1070_33_n_135 | sub_1070_33_n_189));
 assign sub_1070_33_n_196 = ~sub_1070_33_n_195;
 assign sub_1070_33_n_195 = ~sub_1070_33_n_197;
 assign sub_1070_33_n_197 = ~(sub_1070_33_n_176 & (sub_1070_33_n_154 | sub_1070_33_n_189));
 assign T_3_4_ = ((sub_1070_33_n_189 & sub_1070_33_n_136) | ~(sub_1070_33_n_189 | sub_1070_33_n_136));
 assign T_3_3_ = ~((sub_1070_33_n_191 | sub_1070_33_n_113) & ~(sub_1070_33_n_191 & sub_1070_33_n_113));
 assign sub_1070_33_n_192 = ~(sub_1070_33_n_185 | ~sub_1070_33_n_158);
 assign sub_1070_33_n_191 = ~(sub_1070_33_n_66 | (sub_1070_33_n_172 & sub_1070_33_n_83));
 assign sub_1070_33_n_190 = ~(sub_1070_33_n_175 & (sub_1070_33_n_182 | sub_1070_33_n_159));
 assign sub_1070_33_n_189 = ~(sub_1070_33_n_144 | (sub_1070_33_n_172 & sub_1070_33_n_110));
 assign sub_1070_33_n_188 = ~(sub_1070_33_n_186 & ~sub_1070_33_n_32);
 assign T_3_2_ = ~((sub_1070_33_n_172 | sub_1070_33_n_138) & ~(sub_1070_33_n_172 & sub_1070_33_n_138));
 assign sub_1070_33_n_186 = ~(sub_1070_33_n_183 & ~sub_1070_33_n_126);
 assign sub_1070_33_n_185 = ~(sub_1070_33_n_174 | (~sub_1070_33_n_161 & sub_1070_33_n_45));
 assign sub_1070_33_n_184 = ~(sub_1070_33_n_156 & (sub_1070_33_n_177 | sub_1070_33_n_162));
 assign sub_1070_33_n_183 = ~sub_1070_33_n_182;
 assign sub_1070_33_n_182 = ~(sub_1070_33_n_147 | (sub_1070_33_n_166 & sub_1070_33_n_115));
 assign sub_1070_33_n_181 = ~(sub_1070_33_n_167 & sub_1070_33_n_170);
 assign sub_1070_33_n_180 = ~(sub_1070_33_n_168 | ~sub_1070_33_n_127);
 assign sub_1070_33_n_179 = ~(sub_1070_33_n_169 & sub_1070_33_n_158);
 assign sub_1070_33_n_178 = ~sub_1070_33_n_177;
 assign sub_1070_33_n_177 = ~(sub_1070_33_n_148 | (sub_1070_33_n_150 & sub_1070_33_n_120));
 assign sub_1070_33_n_176 = ~(sub_1070_33_n_146 | (sub_1070_33_n_152 & sub_1070_33_n_137));
 assign sub_1070_33_n_175 = ~(sub_1070_33_n_145 | (sub_1070_33_n_32 & sub_1070_33_n_119));
 assign sub_1070_33_n_174 = ~sub_1070_33_n_173;
 assign sub_1070_33_n_173 = ~(sub_1070_33_n_143 | (sub_1070_33_n_149 & sub_1070_33_n_118));
 assign sub_1070_33_n_172 = ~(sub_1070_33_n_84 & (n_1310 | sub_1070_33_n_85));
 assign T_3_1_ = ~((sub_1070_33_n_112 | sub_1070_33_n_165) & ~(sub_1070_33_n_112 & sub_1070_33_n_165));
 assign sub_1070_33_n_170 = ~(sub_1070_33_n_163 | sub_1070_33_n_162);
 assign sub_1070_33_n_169 = ~(sub_1070_33_n_160 | sub_1070_33_n_161);
 assign sub_1070_33_n_168 = ~sub_1070_33_n_167;
 assign sub_1070_33_n_167 = ~(sub_1070_33_n_157 | sub_1070_33_n_159);
 assign sub_1070_33_n_166 = ~(sub_1070_33_n_155 | sub_1070_33_n_38);
 assign sub_1070_33_n_165 = ~n_1310;
 assign sub_1070_33_n_164 = ~sub_1070_33_n_163;
 assign sub_1070_33_n_158 = ~sub_1070_33_n_157;
 assign sub_1070_33_n_156 = ~(sub_1070_33_n_123 & sub_1070_33_n_9);
 assign sub_1070_33_n_155 = ~(sub_1070_33_n_124 & ~sub_1070_33_n_95);
 assign sub_1070_33_n_154 = ~(sub_1070_33_n_135 & sub_1070_33_n_137);
 assign sub_1070_33_n_163 = ~(sub_1070_33_n_127 & sub_1070_33_n_120);
 assign sub_1070_33_n_162 = ~(sub_1070_33_n_123 & sub_1070_33_n_13);
 assign sub_1070_33_n_161 = ~(sub_1070_33_n_114 & sub_1070_33_n_118);
 assign sub_1070_33_n_160 = ~(sub_1070_33_n_130 & sub_1070_33_n_134);
 assign sub_1070_33_n_159 = ~(sub_1070_33_n_125 & sub_1070_33_n_119);
 assign sub_1070_33_n_157 = ~(sub_1070_33_n_122 & sub_1070_33_n_115);
 assign sub_1070_33_n_153 = ~sub_1070_33_n_152;
 assign sub_1070_33_n_148 = ~(sub_1070_33_n_20 & (sub_1070_33_n_3 | sub_1070_33_n_90));
 assign sub_1070_33_n_147 = ~(sub_1070_33_n_10 & (sub_1070_33_n_0 | sub_1070_33_n_68));
 assign sub_1070_33_n_146 = ~(sub_1070_33_n_8 & (sub_1070_33_n_4 | sub_1070_33_n_75));
 assign sub_1070_33_n_145 = ~(sub_1070_33_n_19 & (sub_1070_33_n_12 | sub_1070_33_n_91));
 assign sub_1070_33_n_144 = ~(sub_1070_33_n_106 & (sub_1070_33_n_7 | sub_1070_33_n_69));
 assign sub_1070_33_n_143 = ~(sub_1070_33_n_15 & (sub_1070_33_n_73 | sub_1070_33_n_100));
 assign sub_1070_33_n_152 = ~(sub_1070_33_n_6 & (sub_1070_33_n_1 | sub_1070_33_n_92));
 assign sub_1070_33_n_151 = ~(sub_1070_33_n_105 | (sub_1070_33_n_5 & sub_1070_33_n_18));
 assign sub_1070_33_n_150 = ~(sub_1070_33_n_2 & (sub_1070_33_n_101 | sub_1070_33_n_89));
 assign sub_1070_33_n_149 = ~(sub_1070_33_n_16 & (sub_1070_33_n_11 | sub_1070_33_n_76));
 assign sub_1070_33_n_133 = ~sub_1070_33_n_132;
 assign sub_1070_33_n_126 = ~sub_1070_33_n_125;
 assign sub_1070_33_n_124 = ~(sub_1070_33_n_54 & ~sub_1070_33_n_56);
 assign sub_1070_33_n_142 = ~(sub_1070_33_n_14 & sub_1070_33_n_53);
 assign sub_1070_33_n_141 = ~(sub_1070_33_n_21 & sub_1070_33_n_94);
 assign sub_1070_33_n_140 = ~(sub_1070_33_n_75 | ~sub_1070_33_n_8);
 assign sub_1070_33_n_139 = ~(sub_1070_33_n_68 | ~sub_1070_33_n_10);
 assign sub_1070_33_n_138 = ~(sub_1070_33_n_7 & sub_1070_33_n_83);
 assign sub_1070_33_n_137 = ~(sub_1070_33_n_67 | sub_1070_33_n_75);
 assign sub_1070_33_n_136 = ~(sub_1070_33_n_79 | ~sub_1070_33_n_1);
 assign sub_1070_33_n_135 = ~(sub_1070_33_n_79 | sub_1070_33_n_92);
 assign sub_1070_33_n_134 = ~(sub_1070_33_n_97 | sub_1070_33_n_86);
 assign sub_1070_33_n_132 = ~(sub_1070_33_n_54 & sub_1070_33_n_96);
 assign sub_1070_33_n_131 = ~(sub_1070_33_n_76 | ~sub_1070_33_n_16);
 assign sub_1070_33_n_130 = ~(sub_1070_33_n_72 | sub_1070_33_n_104);
 assign sub_1070_33_n_129 = ~(sub_1070_33_n_70 | sub_1070_33_n_71);
 assign sub_1070_33_n_128 = ~(sub_1070_33_n_17 | sub_1070_33_n_86);
 assign sub_1070_33_n_127 = ~(sub_1070_33_n_98 | ~sub_1070_33_n_88);
 assign sub_1070_33_n_125 = ~(sub_1070_33_n_93 | ~sub_1070_33_n_53);
 assign sub_1070_33_n_110 = ~(sub_1070_33_n_82 | sub_1070_33_n_69);
 assign T_3_0_ = (sub_1070_33_n_65 | (sub_1070_33_n_58 & {in2[3]}));
 assign sub_1070_33_n_123 = ~(n_833 | (n_1276 | n_1364));
 assign sub_1070_33_n_122 = ~(sub_1070_33_n_81 | ~sub_1070_33_n_96);
 assign sub_1070_33_n_121 = ~(sub_1070_33_n_105 | sub_1070_33_n_104);
 assign sub_1070_33_n_120 = ~(sub_1070_33_n_51 | sub_1070_33_n_90);
 assign sub_1070_33_n_119 = ~(sub_1070_33_n_52 | sub_1070_33_n_91);
 assign sub_1070_33_n_118 = ~(sub_1070_33_n_80 | sub_1070_33_n_100);
 assign sub_1070_33_n_117 = ~(sub_1070_33_n_103 | sub_1070_33_n_97);
 assign sub_1070_33_n_116 = ~(sub_1070_33_n_101 & sub_1070_33_n_99);
 assign sub_1070_33_n_115 = ~(sub_1070_33_n_78 | sub_1070_33_n_68);
 assign sub_1070_33_n_114 = ~(sub_1070_33_n_71 | sub_1070_33_n_76);
 assign sub_1070_33_n_113 = ~(sub_1070_33_n_69 | ~sub_1070_33_n_106);
 assign sub_1070_33_n_112 = ~(sub_1070_33_n_84 & (~n_1353 | R_4_0_));
 assign sub_1070_33_n_111 = ~(sub_1070_33_n_74 | sub_1070_33_n_80);
 assign sub_1070_33_n_108 = ~sub_1070_33_n_107;
 assign sub_1070_33_n_104 = ~sub_1070_33_n_18;
 assign sub_1070_33_n_102 = ~sub_1070_33_n_101;
 assign sub_1070_33_n_99 = ~sub_1070_33_n_98;
 assign sub_1070_33_n_96 = ~sub_1070_33_n_95;
 assign sub_1070_33_n_94 = ~sub_1070_33_n_93;
 assign sub_1070_33_n_89 = ~sub_1070_33_n_88;
 assign sub_1070_33_n_87 = ~sub_1070_33_n_4;
 assign sub_1070_33_n_85 = ~(R_4_0_ | ~n_1353);
 assign sub_1070_33_n_107 = ~(sub_1070_33_n_56 & R_4_15_);
 assign sub_1070_33_n_106 = ~(R_4_2_ & ~n_1116);
 assign sub_1070_33_n_105 = ~(n_1165 | sub_1070_33_n_64);
 assign sub_1070_33_n_103 = ~(n_1348 | sub_1070_33_n_63);
 assign sub_1070_33_n_101 = ~(R_4_23_ & ~n_1062);
 assign sub_1070_33_n_100 = ~(R_4_14_ | ~n_1094);
 assign sub_1070_33_n_98 = ~(R_4_23_ | ~n_1062);
 assign sub_1070_33_n_97 = ~(R_4_9_ | ~n_1348);
 assign sub_1070_33_n_54 = ~(R_4_16_ & ~n_1175);
 assign sub_1070_33_n_95 = ~(R_4_16_ | ~n_1175);
 assign sub_1070_33_n_93 = ~(R_4_19_ | ~n_1215);
 assign sub_1070_33_n_92 = ~(R_4_4_ | ~n_1052);
 assign sub_1070_33_n_91 = ~(R_4_22_ | ~n_1295);
 assign sub_1070_33_n_90 = ~(R_4_26_ | ~n_1245);
 assign sub_1070_33_n_88 = ~(sub_1070_33_n_57 & ~sub_1070_33_n_61);
 assign sub_1070_33_n_53 = ~(sub_1070_33_n_62 & ~sub_1070_33_n_59);
 assign sub_1070_33_n_86 = ~(R_4_10_ | ~n_1068);
 assign sub_1070_33_n_83 = ~sub_1070_33_n_82;
 assign sub_1070_33_n_77 = ~sub_1070_33_n_0;
 assign sub_1070_33_n_74 = ~sub_1070_33_n_73;
 assign sub_1070_33_n_70 = ~sub_1070_33_n_11;
 assign sub_1070_33_n_66 = ~sub_1070_33_n_7;
 assign sub_1070_33_n_84 = ~(R_4_0_ & ~n_1353);
 assign sub_1070_33_n_82 = ~(R_4_1_ | ~n_1104);
 assign sub_1070_33_n_81 = ~(R_4_15_ | ~n_1139);
 assign sub_1070_33_n_80 = ~(R_4_13_ | ~n_1185);
 assign sub_1070_33_n_79 = ~(R_4_3_ | ~n_1343);
 assign sub_1070_33_n_78 = ~(R_4_17_ | ~n_1034);
 assign sub_1070_33_n_76 = ~(R_4_12_ | ~n_1262);
 assign sub_1070_33_n_75 = ~(R_4_6_ | ~n_1170);
 assign sub_1070_33_n_52 = ~(R_4_21_ | ~n_1180);
 assign sub_1070_33_n_73 = ~(sub_1070_33_n_60 & R_4_13_);
 assign sub_1070_33_n_72 = ~(R_4_7_ | ~n_1220);
 assign sub_1070_33_n_71 = ~(R_4_11_ | ~n_1029);
 assign sub_1070_33_n_51 = ~(R_4_25_ | ~n_1089);
 assign sub_1070_33_n_69 = ~(R_4_2_ | ~n_1116);
 assign sub_1070_33_n_68 = ~(R_4_18_ | ~n_1305);
 assign sub_1070_33_n_67 = ~(R_4_5_ | ~n_1099);
 assign sub_1070_33_n_65 = ~({in2[3]} | sub_1070_33_n_58);
 assign sub_1070_33_n_64 = ~R_4_8_;
 assign sub_1070_33_n_63 = ~R_4_9_;
 assign sub_1070_33_n_62 = ~R_4_20_;
 assign sub_1070_33_n_61 = ~n_1374;
 assign sub_1070_33_n_60 = ~n_1185;
 assign sub_1070_33_n_59 = ~n_1369;
 assign sub_1070_33_n_58 = ~{in1[0]};
 assign sub_1070_33_n_57 = ~R_4_24_;
 assign sub_1070_33_n_56 = ~n_1139;
 assign sub_1070_33_n_50 = ~(sub_1070_33_n_74 | (~sub_1070_33_n_80 & ~sub_1070_33_n_41));
 assign sub_1070_33_n_49 = ~(sub_1070_33_n_21 & ~(sub_1070_33_n_94 & sub_1070_33_n_214));
 assign sub_1070_33_n_48 = ~(sub_1070_33_n_188 | (~sub_1070_33_n_126 & ~sub_1070_33_n_202));
 assign sub_1070_33_n_47 = (sub_1070_33_n_150 | (sub_1070_33_n_127 & sub_1070_33_n_190));
 assign sub_1070_33_n_46 = ~(sub_1070_33_n_43 & sub_1070_33_n_151);
 assign sub_1070_33_n_45 = ~(sub_1070_33_n_30 & (~sub_1070_33_n_134 | sub_1070_33_n_151));
 assign T_3_15_ = (sub_1070_33_n_50 ^ sub_1070_33_n_40);
 assign sub_1070_33_n_43 = ~(sub_1070_33_n_197 & sub_1070_33_n_130);
 assign sub_1070_33_n_42 = ~(sub_1070_33_n_206 & sub_1070_33_n_122);
 assign sub_1070_33_n_41 = ~(sub_1070_33_n_149 | (sub_1070_33_n_114 & sub_1070_33_n_210));
 assign sub_1070_33_n_40 = ~(sub_1070_33_n_15 & ~sub_1070_33_n_100);
 assign sub_1070_33_n_39 = ~(sub_1070_33_n_103 | (~sub_1070_33_n_97 & sub_1070_33_n_46));
 assign sub_1070_33_n_38 = ~(R_4_15_ | ~sub_1070_33_n_54);
 assign sub_1070_33_n_37 = ~(sub_1070_33_n_6 & ~sub_1070_33_n_92);
 assign sub_1070_33_n_36 = (sub_1070_33_n_5 | sub_1070_33_n_72);
 assign sub_1070_33_n_35 = ~(sub_1070_33_n_52 | ~sub_1070_33_n_12);
 assign sub_1070_33_n_34 = ~(sub_1070_33_n_19 & ~sub_1070_33_n_91);
 assign sub_1070_33_n_33 = ~(sub_1070_33_n_20 & ~sub_1070_33_n_90);
 assign sub_1070_33_n_32 = ~(sub_1070_33_n_14 & (~sub_1070_33_n_53 | sub_1070_33_n_21));
 assign sub_1070_33_n_31 = ~(sub_1070_33_n_51 | ~sub_1070_33_n_3);
 assign sub_1070_33_n_30 = ~(sub_1070_33_n_17 | (~sub_1070_33_n_86 & sub_1070_33_n_103));
 assign sub_1070_33_n_29 = ~(sub_1070_33_n_89 | ~sub_1070_33_n_2);
 assign sub_1070_33_n_28 = ~(sub_1070_33_n_9 | ~sub_1070_33_n_13);
 assign sub_1070_33_n_27 = ~(sub_1070_33_n_107 & ~sub_1070_33_n_81);
 assign sub_1070_33_n_26 = ~(sub_1070_33_n_1 & (sub_1070_33_n_79 | sub_1070_33_n_189));
 assign sub_1070_33_n_25 = ~(sub_1070_33_n_0 & ~sub_1070_33_n_78);
 assign sub_1070_33_n_24 = ~(sub_1070_33_n_12 & (sub_1070_33_n_52 | sub_1070_33_n_48));
 assign sub_1070_33_n_23 = ~(sub_1070_33_n_3 & (sub_1070_33_n_51 | sub_1070_33_n_220));
 assign sub_1070_33_n_22 = ~(sub_1070_33_n_4 & ~sub_1070_33_n_67);
 assign sub_1070_33_n_21 = ~(R_4_19_ & ~n_1215);
 assign sub_1070_33_n_20 = ~(R_4_26_ & ~n_1245);
 assign sub_1070_33_n_19 = ~(R_4_22_ & ~n_1295);
 assign sub_1070_33_n_18 = ~(sub_1070_33_n_64 & n_1165);
 assign sub_1070_33_n_17 = ~(n_1068 | ~R_4_10_);
 assign sub_1070_33_n_16 = ~(R_4_12_ & ~n_1262);
 assign sub_1070_33_n_15 = ~(R_4_14_ & ~n_1094);
 assign sub_1070_33_n_14 = ~(sub_1070_33_n_59 & ~sub_1070_33_n_62);
 assign sub_1070_33_n_13 = ~(n_1300 & ~R_4_27_);
 assign sub_1070_33_n_12 = ~(R_4_21_ & ~n_1180);
 assign sub_1070_33_n_11 = ~(R_4_11_ & ~n_1029);
 assign sub_1070_33_n_10 = ~(R_4_18_ & ~n_1305);
 assign sub_1070_33_n_9 = ~(n_1300 | ~R_4_27_);
 assign sub_1070_33_n_8 = ~(R_4_6_ & ~n_1170);
 assign sub_1070_33_n_7 = ~(R_4_1_ & ~n_1104);
 assign sub_1070_33_n_6 = ~(R_4_4_ & ~n_1052);
 assign sub_1070_33_n_5 = ~(n_1220 | ~R_4_7_);
 assign sub_1070_33_n_4 = ~(R_4_5_ & ~n_1099);
 assign sub_1070_33_n_3 = ~(R_4_25_ & ~n_1089);
 assign sub_1070_33_n_2 = ~(sub_1070_33_n_61 & ~sub_1070_33_n_57);
 assign sub_1070_33_n_1 = ~(R_4_3_ & ~n_1343);
 assign sub_1070_33_n_0 = ~(R_4_17_ & ~n_1034);
 assign T_2_23_ = ~(sub_1100_32_n_260 & sub_1100_32_n_37);
 assign T_2_29_ = ((sub_1100_32_n_262 & sub_1100_32_n_27) | ~(sub_1100_32_n_262 | sub_1100_32_n_27));
 assign T_2_27_ = ((sub_1100_32_n_261 & sub_1100_32_n_28) | ~(sub_1100_32_n_261 | sub_1100_32_n_28));
 assign sub_1100_32_n_262 = ~(sub_1100_32_n_79 | (sub_1100_32_n_32 & sub_1100_32_n_67));
 assign sub_1100_32_n_261 = ~(sub_1100_32_n_75 | (sub_1100_32_n_249 & sub_1100_32_n_82));
 assign sub_1100_32_n_260 = ~(sub_1100_32_n_252 & ~sub_1100_32_n_178);
 assign T_2_22_ = ((sub_1100_32_n_248 & sub_1100_32_n_19) | ~(sub_1100_32_n_248 | sub_1100_32_n_19));
 assign T_2_21_ = ((sub_1100_32_n_250 & sub_1100_32_n_163) | ~(sub_1100_32_n_250 | sub_1100_32_n_163));
 assign T_2_19_ = ((sub_1100_32_n_251 & sub_1100_32_n_23) | ~(sub_1100_32_n_251 | sub_1100_32_n_23));
 assign T_2_15_ = ((sub_1100_32_n_36 & sub_1100_32_n_153) | ~(sub_1100_32_n_36 | sub_1100_32_n_153));
 assign T_2_28_ = ((sub_1100_32_n_32 & sub_1100_32_n_142) | ~(sub_1100_32_n_32 | sub_1100_32_n_142));
 assign T_2_26_ = ((sub_1100_32_n_249 & sub_1100_32_n_138) | ~(sub_1100_32_n_249 | sub_1100_32_n_138));
 assign T_2_25_ = ~((sub_1100_32_n_35 | sub_1100_32_n_135) & ~(sub_1100_32_n_35 & sub_1100_32_n_135));
 assign sub_1100_32_n_252 = ~(sub_1100_32_n_248 & ~sub_1100_32_n_71);
 assign sub_1100_32_n_251 = ~(sub_1100_32_n_5 & (~sub_1100_32_n_0 | sub_1100_32_n_30));
 assign sub_1100_32_n_250 = ~(sub_1100_32_n_43 & (~sub_1100_32_n_104 | sub_1100_32_n_235));
 assign sub_1100_32_n_249 = ~(sub_1100_32_n_181 & (~sub_1100_32_n_144 | sub_1100_32_n_234));
 assign sub_1100_32_n_248 = ~(sub_1100_32_n_175 & (~sub_1100_32_n_154 | sub_1100_32_n_235));
 assign T_2_24_ = ~((sub_1100_32_n_234 | sub_1100_32_n_134) & ~(sub_1100_32_n_234 & sub_1100_32_n_134));
 assign T_2_18_ = ~((sub_1100_32_n_30 | sub_1100_32_n_160) & ~(sub_1100_32_n_30 & sub_1100_32_n_160));
 assign T_2_17_ = ~((sub_1100_32_n_34 | sub_1100_32_n_157) & ~(sub_1100_32_n_34 & sub_1100_32_n_157));
 assign T_2_14_ = ~((sub_1100_32_n_237 | sub_1100_32_n_151) & ~(sub_1100_32_n_237 & sub_1100_32_n_151));
 assign T_2_13_ = ~((sub_1100_32_n_239 | sub_1100_32_n_152) & ~(sub_1100_32_n_239 & sub_1100_32_n_152));
 assign T_2_11_ = ((sub_1100_32_n_238 & sub_1100_32_n_150) | ~(sub_1100_32_n_238 | sub_1100_32_n_150));
 assign T_2_20_ = ((sub_1100_32_n_235 & sub_1100_32_n_22) | ~(sub_1100_32_n_235 | sub_1100_32_n_22));
 assign T_2_32_ = ~sub_1100_32_n_236;
 assign sub_1100_32_n_236 = ~(sub_1100_32_n_226 & sub_1100_32_n_207);
 assign sub_1100_32_n_239 = ~(sub_1100_32_n_125 | (~sub_1100_32_n_102 & sub_1100_32_n_224));
 assign sub_1100_32_n_238 = ~(sub_1100_32_n_123 | (~sub_1100_32_n_117 & sub_1100_32_n_222));
 assign sub_1100_32_n_237 = ~(sub_1100_32_n_173 | (~sub_1100_32_n_24 & sub_1100_32_n_224));
 assign T_2_16_ = ((sub_1100_32_n_44 & sub_1100_32_n_156) | ~(sub_1100_32_n_44 | sub_1100_32_n_156));
 assign T_2_7_ = ((sub_1100_32_n_220 & sub_1100_32_n_25) | ~(sub_1100_32_n_220 | sub_1100_32_n_25));
 assign T_2_12_ = ((sub_1100_32_n_225 & sub_1100_32_n_161) | ~(sub_1100_32_n_225 | sub_1100_32_n_161));
 assign T_2_10_ = ((sub_1100_32_n_223 & sub_1100_32_n_147) | ~(sub_1100_32_n_223 | sub_1100_32_n_147));
 assign T_2_9_ = ((sub_1100_32_n_221 & sub_1100_32_n_26) | ~(sub_1100_32_n_221 | sub_1100_32_n_26));
 assign sub_1100_32_n_235 = ~(sub_1100_32_n_227 | ~sub_1100_32_n_197);
 assign sub_1100_32_n_234 = ~(sub_1100_32_n_203 | (~sub_1100_32_n_190 & sub_1100_32_n_219));
 assign sub_1100_32_n_228 = ~(sub_1100_32_n_44 | ~sub_1100_32_n_143);
 assign sub_1100_32_n_227 = ~(sub_1100_32_n_44 | ~sub_1100_32_n_185);
 assign sub_1100_32_n_226 = ~(sub_1100_32_n_219 & ~sub_1100_32_n_200);
 assign sub_1100_32_n_225 = ~sub_1100_32_n_224;
 assign sub_1100_32_n_224 = ~(sub_1100_32_n_33 & ~sub_1100_32_n_39);
 assign sub_1100_32_n_223 = ~sub_1100_32_n_222;
 assign sub_1100_32_n_222 = ~(sub_1100_32_n_215 & ~sub_1100_32_n_172);
 assign sub_1100_32_n_221 = ~(sub_1100_32_n_69 | (~sub_1100_32_n_116 & sub_1100_32_n_213));
 assign sub_1100_32_n_220 = ~(sub_1100_32_n_11 & (~sub_1100_32_n_85 | sub_1100_32_n_29));
 assign sub_1100_32_n_44 = ~sub_1100_32_n_219;
 assign sub_1100_32_n_219 = ~(sub_1100_32_n_31 & sub_1100_32_n_214);
 assign T_2_6_ = ((sub_1100_32_n_29 & sub_1100_32_n_130) | ~(sub_1100_32_n_29 | sub_1100_32_n_130));
 assign T_2_5_ = ~((sub_1100_32_n_212 | sub_1100_32_n_155) & ~(sub_1100_32_n_212 & sub_1100_32_n_155));
 assign T_2_8_ = ~((sub_1100_32_n_213 | sub_1100_32_n_149) & ~(sub_1100_32_n_213 & sub_1100_32_n_149));
 assign sub_1100_32_n_215 = ~(sub_1100_32_n_213 & ~sub_1100_32_n_132);
 assign sub_1100_32_n_214 = ~(sub_1100_32_n_213 & ~sub_1100_32_n_191);
 assign sub_1100_32_n_213 = ~(sub_1100_32_n_196 & (sub_1100_32_n_179 | sub_1100_32_n_205));
 assign sub_1100_32_n_212 = ~(sub_1100_32_n_209 | ~sub_1100_32_n_122);
 assign T_2_4_ = ((sub_1100_32_n_205 & sub_1100_32_n_141) | ~(sub_1100_32_n_205 | sub_1100_32_n_141));
 assign T_2_3_ = ~((sub_1100_32_n_206 | sub_1100_32_n_162) & ~(sub_1100_32_n_206 & sub_1100_32_n_162));
 assign sub_1100_32_n_209 = ~(sub_1100_32_n_205 | ~sub_1100_32_n_114);
 assign sub_1100_32_n_208 = ~(sub_1100_32_n_205 | ~sub_1100_32_n_140);
 assign sub_1100_32_n_207 = ~(sub_1100_32_n_202 | (sub_1100_32_n_203 & sub_1100_32_n_193));
 assign sub_1100_32_n_206 = ~(sub_1100_32_n_91 | (~sub_1100_32_n_90 & sub_1100_32_n_201));
 assign sub_1100_32_n_205 = ~(sub_1100_32_n_169 | (sub_1100_32_n_128 & sub_1100_32_n_201));
 assign T_2_2_ = ~((sub_1100_32_n_201 | sub_1100_32_n_20) & ~(sub_1100_32_n_201 & sub_1100_32_n_20));
 assign sub_1100_32_n_203 = ~(sub_1100_32_n_194 & (sub_1100_32_n_197 | sub_1100_32_n_183));
 assign sub_1100_32_n_202 = ((sub_1100_32_n_170 & sub_1100_32_n_94) | ~(sub_1100_32_n_195 | sub_1100_32_n_21));
 assign sub_1100_32_n_201 = ~(sub_1100_32_n_198 & sub_1100_32_n_93);
 assign sub_1100_32_n_200 = ~(sub_1100_32_n_189 & sub_1100_32_n_193);
 assign T_2_1_ = ((sub_1100_32_n_129 & n_1255) | ~(sub_1100_32_n_129 | n_1255));
 assign sub_1100_32_n_198 = ~(sub_1100_32_n_192 | (n_1255 & R_3_0_));
 assign sub_1100_32_n_197 = ~(sub_1100_32_n_168 | (~sub_1100_32_n_145 & sub_1100_32_n_182));
 assign sub_1100_32_n_196 = ~(sub_1100_32_n_166 | (sub_1100_32_n_176 & sub_1100_32_n_139));
 assign sub_1100_32_n_195 = ~(sub_1100_32_n_167 | (sub_1100_32_n_180 & sub_1100_32_n_164));
 assign sub_1100_32_n_194 = ~(sub_1100_32_n_171 | (sub_1100_32_n_131 & sub_1100_32_n_174));
 assign sub_1100_32_n_193 = ~(sub_1100_32_n_21 | sub_1100_32_n_187);
 assign sub_1100_32_n_192 = ~(n_1353 | ~n_1255);
 assign sub_1100_32_n_191 = ~(sub_1100_32_n_188 & sub_1100_32_n_186);
 assign sub_1100_32_n_190 = ~sub_1100_32_n_189;
 assign sub_1100_32_n_189 = ~(sub_1100_32_n_184 | sub_1100_32_n_183);
 assign sub_1100_32_n_185 = ~sub_1100_32_n_184;
 assign sub_1100_32_n_181 = ~sub_1100_32_n_180;
 assign sub_1100_32_n_179 = ~(sub_1100_32_n_140 & sub_1100_32_n_139);
 assign sub_1100_32_n_178 = ~(sub_1100_32_n_133 & sub_1100_32_n_97);
 assign sub_1100_32_n_177 = ~(sub_1100_32_n_95 & (sub_1100_32_n_8 | sub_1100_32_n_106));
 assign sub_1100_32_n_188 = ~(sub_1100_32_n_132 | sub_1100_32_n_158);
 assign sub_1100_32_n_187 = ~(sub_1100_32_n_144 & sub_1100_32_n_164);
 assign sub_1100_32_n_186 = ~(sub_1100_32_n_24 | sub_1100_32_n_136);
 assign sub_1100_32_n_184 = ~(sub_1100_32_n_143 & sub_1100_32_n_146);
 assign sub_1100_32_n_183 = ~(sub_1100_32_n_154 & sub_1100_32_n_131);
 assign sub_1100_32_n_182 = ~(sub_1100_32_n_4 & (sub_1100_32_n_76 | sub_1100_32_n_88));
 assign sub_1100_32_n_180 = ~(sub_1100_32_n_10 & (sub_1100_32_n_107 | sub_1100_32_n_120));
 assign sub_1100_32_n_175 = ~sub_1100_32_n_174;
 assign sub_1100_32_n_171 = ~(sub_1100_32_n_2 & (sub_1100_32_n_97 | sub_1100_32_n_65));
 assign sub_1100_32_n_170 = ~(sub_1100_32_n_12 & (sub_1100_32_n_78 | sub_1100_32_n_86));
 assign sub_1100_32_n_169 = ~(sub_1100_32_n_1 & (sub_1100_32_n_42 | sub_1100_32_n_98));
 assign sub_1100_32_n_168 = ~(sub_1100_32_n_18 & (sub_1100_32_n_5 | sub_1100_32_n_112));
 assign sub_1100_32_n_167 = ~(sub_1100_32_n_9 & (sub_1100_32_n_74 | sub_1100_32_n_83));
 assign sub_1100_32_n_166 = ~(sub_1100_32_n_14 & (sub_1100_32_n_11 | sub_1100_32_n_121));
 assign sub_1100_32_n_165 = ~(sub_1100_32_n_92 & (sub_1100_32_n_7 | sub_1100_32_n_100));
 assign sub_1100_32_n_176 = ~(sub_1100_32_n_15 & (sub_1100_32_n_122 | sub_1100_32_n_110));
 assign sub_1100_32_n_174 = ~(sub_1100_32_n_3 & (sub_1100_32_n_43 | sub_1100_32_n_68));
 assign sub_1100_32_n_173 = ~(sub_1100_32_n_17 & (sub_1100_32_n_124 | sub_1100_32_n_118));
 assign sub_1100_32_n_172 = ~(sub_1100_32_n_126 & (sub_1100_32_n_41 | sub_1100_32_n_109));
 assign sub_1100_32_n_159 = ~sub_1100_32_n_158;
 assign sub_1100_32_n_148 = ~(sub_1100_32_n_66 | sub_1100_32_n_86);
 assign sub_1100_32_n_164 = ~(sub_1100_32_n_81 | sub_1100_32_n_83);
 assign sub_1100_32_n_163 = ~(sub_1100_32_n_3 & sub_1100_32_n_40);
 assign sub_1100_32_n_162 = ~(sub_1100_32_n_98 | ~sub_1100_32_n_1);
 assign sub_1100_32_n_161 = ~(sub_1100_32_n_125 | sub_1100_32_n_102);
 assign sub_1100_32_n_160 = (sub_1100_32_n_5 & sub_1100_32_n_0);
 assign sub_1100_32_n_158 = ~(sub_1100_32_n_13 & sub_1100_32_n_105);
 assign sub_1100_32_n_157 = ~(sub_1100_32_n_88 | ~sub_1100_32_n_4);
 assign sub_1100_32_n_156 = ~(sub_1100_32_n_77 | sub_1100_32_n_89);
 assign sub_1100_32_n_155 = ~(sub_1100_32_n_110 | ~sub_1100_32_n_15);
 assign sub_1100_32_n_154 = ~(sub_1100_32_n_103 | ~sub_1100_32_n_40);
 assign sub_1100_32_n_153 = ~(sub_1100_32_n_100 | ~sub_1100_32_n_92);
 assign sub_1100_32_n_152 = ~(sub_1100_32_n_118 | ~sub_1100_32_n_17);
 assign sub_1100_32_n_151 = ~(sub_1100_32_n_80 | sub_1100_32_n_73);
 assign sub_1100_32_n_150 = ~(sub_1100_32_n_106 | ~sub_1100_32_n_95);
 assign sub_1100_32_n_149 = ~(sub_1100_32_n_41 & sub_1100_32_n_115);
 assign sub_1100_32_n_146 = ~sub_1100_32_n_145;
 assign sub_1100_32_n_137 = ~sub_1100_32_n_136;
 assign sub_1100_32_n_128 = ~(sub_1100_32_n_90 | sub_1100_32_n_98);
 assign T_2_0_ = ~(sub_1100_32_n_96 & (~{in2[2]} | {in1[0]}));
 assign sub_1100_32_n_147 = ~(sub_1100_32_n_123 | sub_1100_32_n_117);
 assign sub_1100_32_n_145 = ~(sub_1100_32_n_0 & sub_1100_32_n_111);
 assign sub_1100_32_n_144 = ~(sub_1100_32_n_70 | ~sub_1100_32_n_119);
 assign sub_1100_32_n_143 = ~(sub_1100_32_n_89 | ~sub_1100_32_n_87);
 assign sub_1100_32_n_142 = ~(sub_1100_32_n_78 & sub_1100_32_n_67);
 assign sub_1100_32_n_141 = (sub_1100_32_n_122 & sub_1100_32_n_114);
 assign sub_1100_32_n_140 = ~(sub_1100_32_n_113 | sub_1100_32_n_110);
 assign sub_1100_32_n_139 = ~(sub_1100_32_n_84 | sub_1100_32_n_121);
 assign sub_1100_32_n_138 = ~(sub_1100_32_n_74 & sub_1100_32_n_82);
 assign sub_1100_32_n_136 = ~(sub_1100_32_n_72 & sub_1100_32_n_99);
 assign sub_1100_32_n_135 = ~(sub_1100_32_n_120 | ~sub_1100_32_n_10);
 assign sub_1100_32_n_134 = ~(sub_1100_32_n_108 | sub_1100_32_n_70);
 assign sub_1100_32_n_133 = ~(sub_1100_32_n_65 | ~sub_1100_32_n_2);
 assign sub_1100_32_n_132 = ~(sub_1100_32_n_115 & sub_1100_32_n_6);
 assign sub_1100_32_n_131 = ~(sub_1100_32_n_71 | sub_1100_32_n_65);
 assign sub_1100_32_n_130 = (sub_1100_32_n_11 & sub_1100_32_n_85);
 assign sub_1100_32_n_129 = ~(sub_1100_32_n_93 & (~n_1353 | R_3_0_));
 assign sub_1100_32_n_125 = ~sub_1100_32_n_124;
 assign sub_1100_32_n_123 = ~sub_1100_32_n_8;
 assign sub_1100_32_n_120 = ~sub_1100_32_n_119;
 assign sub_1100_32_n_117 = ~sub_1100_32_n_13;
 assign sub_1100_32_n_116 = ~sub_1100_32_n_115;
 assign sub_1100_32_n_114 = ~sub_1100_32_n_113;
 assign sub_1100_32_n_112 = ~sub_1100_32_n_111;
 assign sub_1100_32_n_108 = ~sub_1100_32_n_107;
 assign sub_1100_32_n_106 = ~sub_1100_32_n_105;
 assign sub_1100_32_n_104 = ~sub_1100_32_n_103;
 assign sub_1100_32_n_102 = ~sub_1100_32_n_16;
 assign sub_1100_32_n_101 = ~sub_1100_32_n_43;
 assign sub_1100_32_n_100 = ~sub_1100_32_n_99;
 assign sub_1100_32_n_126 = ~(sub_1100_32_n_55 & R_3_8_);
 assign sub_1100_32_n_124 = ~(R_3_11_ & ~n_1029);
 assign sub_1100_32_n_122 = ~(R_3_3_ & ~n_1343);
 assign sub_1100_32_n_121 = ~(R_3_6_ | ~n_1170);
 assign sub_1100_32_n_119 = ~(sub_1100_32_n_59 & ~sub_1100_32_n_47);
 assign sub_1100_32_n_118 = ~(R_3_12_ | ~n_1262);
 assign sub_1100_32_n_115 = ~(sub_1100_32_n_61 & ~sub_1100_32_n_57);
 assign sub_1100_32_n_113 = ~(R_3_3_ | ~n_1343);
 assign sub_1100_32_n_111 = ~(sub_1100_32_n_64 & ~sub_1100_32_n_48);
 assign sub_1100_32_n_110 = ~(R_3_4_ | ~n_1052);
 assign sub_1100_32_n_109 = ~(R_3_8_ | ~n_1165);
 assign sub_1100_32_n_107 = ~(R_3_23_ & ~n_1062);
 assign sub_1100_32_n_105 = ~(sub_1100_32_n_62 & ~sub_1100_32_n_50);
 assign sub_1100_32_n_103 = ~(R_3_19_ | ~n_1215);
 assign sub_1100_32_n_99 = ~(sub_1100_32_n_46 & ~sub_1100_32_n_63);
 assign sub_1100_32_n_98 = ~(R_3_2_ | ~n_1116);
 assign sub_1100_32_n_97 = ~(R_3_21_ & ~n_1180);
 assign sub_1100_32_n_96 = ~({in1[0]} & ~{in2[2]});
 assign sub_1100_32_n_91 = ~sub_1100_32_n_42;
 assign sub_1100_32_n_88 = ~sub_1100_32_n_87;
 assign sub_1100_32_n_85 = ~sub_1100_32_n_84;
 assign sub_1100_32_n_82 = ~sub_1100_32_n_81;
 assign sub_1100_32_n_80 = ~sub_1100_32_n_7;
 assign sub_1100_32_n_79 = ~sub_1100_32_n_78;
 assign sub_1100_32_n_77 = ~sub_1100_32_n_76;
 assign sub_1100_32_n_75 = ~sub_1100_32_n_74;
 assign sub_1100_32_n_73 = ~sub_1100_32_n_72;
 assign sub_1100_32_n_69 = ~sub_1100_32_n_41;
 assign sub_1100_32_n_68 = ~sub_1100_32_n_40;
 assign sub_1100_32_n_67 = ~sub_1100_32_n_66;
 assign sub_1100_32_n_95 = ~(sub_1100_32_n_50 & R_3_10_);
 assign sub_1100_32_n_94 = ~(n_833 | n_1276);
 assign sub_1100_32_n_93 = ~(R_3_0_ & ~n_1353);
 assign sub_1100_32_n_92 = ~(sub_1100_32_n_63 & R_3_14_);
 assign sub_1100_32_n_42 = ~(R_3_1_ & ~n_1104);
 assign sub_1100_32_n_90 = ~(R_3_1_ | ~n_1104);
 assign sub_1100_32_n_89 = ~(R_3_15_ | ~n_1139);
 assign sub_1100_32_n_87 = ~(sub_1100_32_n_51 & ~sub_1100_32_n_60);
 assign sub_1100_32_n_86 = ~(R_3_28_ | ~n_1364);
 assign sub_1100_32_n_84 = ~(R_3_5_ | ~n_1099);
 assign sub_1100_32_n_83 = ~(R_3_26_ | ~n_1245);
 assign sub_1100_32_n_81 = ~(R_3_25_ | ~n_1089);
 assign sub_1100_32_n_78 = ~(R_3_27_ & ~n_1300);
 assign sub_1100_32_n_76 = ~(R_3_15_ & ~n_1139);
 assign sub_1100_32_n_74 = ~(R_3_25_ & ~n_1089);
 assign sub_1100_32_n_72 = ~(sub_1100_32_n_53 & ~sub_1100_32_n_58);
 assign sub_1100_32_n_71 = ~(R_3_21_ | ~n_1180);
 assign sub_1100_32_n_70 = ~(R_3_23_ | ~n_1062);
 assign sub_1100_32_n_41 = ~(sub_1100_32_n_57 & R_3_7_);
 assign sub_1100_32_n_40 = ~(sub_1100_32_n_49 & ~sub_1100_32_n_54);
 assign sub_1100_32_n_66 = ~(R_3_27_ | ~n_1300);
 assign sub_1100_32_n_65 = ~(R_3_22_ | ~n_1295);
 assign sub_1100_32_n_64 = ~R_3_18_;
 assign sub_1100_32_n_63 = ~n_1094;
 assign sub_1100_32_n_62 = ~R_3_10_;
 assign sub_1100_32_n_61 = ~R_3_7_;
 assign sub_1100_32_n_60 = ~n_1175;
 assign sub_1100_32_n_59 = ~R_3_24_;
 assign sub_1100_32_n_58 = ~n_1185;
 assign sub_1100_32_n_57 = ~n_1220;
 assign sub_1100_32_n_56 = ~R_3_9_;
 assign sub_1100_32_n_55 = ~n_1165;
 assign sub_1100_32_n_54 = ~n_1369;
 assign sub_1100_32_n_53 = ~R_3_13_;
 assign sub_1100_32_n_52 = ~R_3_17_;
 assign sub_1100_32_n_51 = ~R_3_16_;
 assign sub_1100_32_n_50 = ~n_1068;
 assign sub_1100_32_n_49 = ~R_3_20_;
 assign sub_1100_32_n_48 = ~n_1305;
 assign sub_1100_32_n_47 = ~n_1374;
 assign sub_1100_32_n_46 = ~R_3_14_;
 assign sub_1100_32_n_39 = (sub_1100_32_n_177 | (sub_1100_32_n_172 & sub_1100_32_n_159));
 assign sub_1100_32_n_38 = (sub_1100_32_n_165 | (sub_1100_32_n_173 & sub_1100_32_n_137));
 assign sub_1100_32_n_37 = (sub_1100_32_n_133 | (sub_1100_32_n_97 & sub_1100_32_n_252));
 assign sub_1100_32_n_36 = ~(sub_1100_32_n_80 | (~sub_1100_32_n_73 & ~sub_1100_32_n_237));
 assign sub_1100_32_n_35 = ~(sub_1100_32_n_108 | (~sub_1100_32_n_70 & ~sub_1100_32_n_234));
 assign sub_1100_32_n_34 = ~(sub_1100_32_n_77 | (~sub_1100_32_n_89 & ~sub_1100_32_n_44));
 assign sub_1100_32_n_33 = ~(sub_1100_32_n_213 & sub_1100_32_n_188);
 assign sub_1100_32_n_32 = ~(sub_1100_32_n_195 & (sub_1100_32_n_187 | sub_1100_32_n_234));
 assign sub_1100_32_n_31 = ~(sub_1100_32_n_38 | (sub_1100_32_n_186 & sub_1100_32_n_39));
 assign sub_1100_32_n_30 = ~(sub_1100_32_n_228 | sub_1100_32_n_182);
 assign sub_1100_32_n_29 = ~(sub_1100_32_n_208 | sub_1100_32_n_176);
 assign sub_1100_32_n_28 = ~(sub_1100_32_n_83 | ~sub_1100_32_n_9);
 assign sub_1100_32_n_27 = ~(sub_1100_32_n_86 | ~sub_1100_32_n_12);
 assign sub_1100_32_n_26 = ~(sub_1100_32_n_109 | ~sub_1100_32_n_126);
 assign sub_1100_32_n_25 = ~(sub_1100_32_n_14 & ~sub_1100_32_n_121);
 assign sub_1100_32_n_24 = ~(sub_1100_32_n_16 & ~sub_1100_32_n_118);
 assign sub_1100_32_n_23 = ~(sub_1100_32_n_18 & ~sub_1100_32_n_112);
 assign sub_1100_32_n_22 = ~(sub_1100_32_n_101 | ~sub_1100_32_n_104);
 assign sub_1100_32_n_21 = ~(sub_1100_32_n_148 & sub_1100_32_n_94);
 assign sub_1100_32_n_20 = ~(sub_1100_32_n_42 & ~sub_1100_32_n_90);
 assign sub_1100_32_n_19 = ~(sub_1100_32_n_97 & ~sub_1100_32_n_71);
 assign sub_1100_32_n_18 = ~(sub_1100_32_n_48 & ~sub_1100_32_n_64);
 assign sub_1100_32_n_17 = ~(R_3_12_ & ~n_1262);
 assign sub_1100_32_n_16 = ~(n_1029 & ~R_3_11_);
 assign sub_1100_32_n_43 = ~(R_3_19_ & ~n_1215);
 assign sub_1100_32_n_15 = ~(R_3_4_ & ~n_1052);
 assign sub_1100_32_n_14 = ~(R_3_6_ & ~n_1170);
 assign sub_1100_32_n_13 = ~(sub_1100_32_n_56 & n_1348);
 assign sub_1100_32_n_12 = ~(R_3_28_ & ~n_1364);
 assign sub_1100_32_n_11 = ~(R_3_5_ & ~n_1099);
 assign sub_1100_32_n_10 = ~(sub_1100_32_n_47 & ~sub_1100_32_n_59);
 assign sub_1100_32_n_9 = ~(R_3_26_ & ~n_1245);
 assign sub_1100_32_n_8 = (sub_1100_32_n_56 | n_1348);
 assign sub_1100_32_n_7 = ~(sub_1100_32_n_58 & ~sub_1100_32_n_53);
 assign sub_1100_32_n_6 = (R_3_8_ | sub_1100_32_n_55);
 assign sub_1100_32_n_5 = (sub_1100_32_n_52 | n_1034);
 assign sub_1100_32_n_4 = ~(sub_1100_32_n_60 & ~sub_1100_32_n_51);
 assign sub_1100_32_n_3 = ~(sub_1100_32_n_54 & ~sub_1100_32_n_49);
 assign sub_1100_32_n_2 = ~(R_3_22_ & ~n_1295);
 assign sub_1100_32_n_1 = ~(R_3_2_ & ~n_1116);
 assign sub_1100_32_n_0 = ~(sub_1100_32_n_52 & n_1034);
 assign T_1_30_ = ~(sub_1130_31_n_248 & sub_1130_31_n_250);
 assign T_1_23_ = ~(sub_1130_31_n_247 & sub_1130_31_n_42);
 assign T_1_29_ = ((sub_1130_31_n_19 & sub_1130_31_n_127) | ~(sub_1130_31_n_19 | sub_1130_31_n_127));
 assign T_1_27_ = ~((sub_1130_31_n_249 | sub_1130_31_n_119) & ~(sub_1130_31_n_249 & sub_1130_31_n_119));
 assign sub_1130_31_n_250 = ~(sub_1130_31_n_123 & (~sub_1130_31_n_148 | sub_1130_31_n_237));
 assign sub_1130_31_n_248 = ~(sub_1130_31_n_238 & ~sub_1130_31_n_167);
 assign sub_1130_31_n_247 = ~(sub_1130_31_n_239 & ~sub_1130_31_n_155);
 assign T_1_22_ = ((sub_1130_31_n_233 & sub_1130_31_n_30) | ~(sub_1130_31_n_233 | sub_1130_31_n_30));
 assign sub_1130_31_n_249 = ~(sub_1130_31_n_89 & (~sub_1130_31_n_15 | sub_1130_31_n_34));
 assign T_1_21_ = ((sub_1130_31_n_236 & sub_1130_31_n_23) | ~(sub_1130_31_n_236 | sub_1130_31_n_23));
 assign T_1_19_ = ~((sub_1130_31_n_235 | sub_1130_31_n_17) & ~(sub_1130_31_n_235 & sub_1130_31_n_17));
 assign T_1_15_ = ((sub_1130_31_n_234 & sub_1130_31_n_133) | ~(sub_1130_31_n_234 | sub_1130_31_n_133));
 assign T_1_28_ = ((sub_1130_31_n_232 & sub_1130_31_n_31) | ~(sub_1130_31_n_232 | sub_1130_31_n_31));
 assign T_1_26_ = ((sub_1130_31_n_34 & sub_1130_31_n_25) | ~(sub_1130_31_n_34 | sub_1130_31_n_25));
 assign T_1_25_ = ((sub_1130_31_n_41 & sub_1130_31_n_115) | ~(sub_1130_31_n_41 | sub_1130_31_n_115));
 assign sub_1130_31_n_239 = ~(sub_1130_31_n_233 & ~sub_1130_31_n_97);
 assign sub_1130_31_n_238 = ~sub_1130_31_n_237;
 assign sub_1130_31_n_237 = ~(sub_1130_31_n_232 | ~sub_1130_31_n_126);
 assign sub_1130_31_n_236 = ~(sub_1130_31_n_101 & (~sub_1130_31_n_60 | sub_1130_31_n_222));
 assign sub_1130_31_n_235 = ~(sub_1130_31_n_98 & (~sub_1130_31_n_85 | sub_1130_31_n_224));
 assign sub_1130_31_n_234 = ~(sub_1130_31_n_62 | (sub_1130_31_n_223 & sub_1130_31_n_65));
 assign sub_1130_31_n_233 = ~(sub_1130_31_n_36 & ~sub_1130_31_n_160);
 assign sub_1130_31_n_232 = ~(sub_1130_31_n_177 | (sub_1130_31_n_219 & sub_1130_31_n_163));
 assign T_1_24_ = ((sub_1130_31_n_219 & sub_1130_31_n_114) | ~(sub_1130_31_n_219 | sub_1130_31_n_114));
 assign T_1_18_ = ((sub_1130_31_n_224 & sub_1130_31_n_135) | ~(sub_1130_31_n_224 | sub_1130_31_n_135));
 assign T_1_17_ = ~((sub_1130_31_n_40 | sub_1130_31_n_20) & ~(sub_1130_31_n_40 & sub_1130_31_n_20));
 assign T_1_14_ = ~((sub_1130_31_n_223 | sub_1130_31_n_131) & ~(sub_1130_31_n_223 & sub_1130_31_n_131));
 assign T_1_13_ = ((sub_1130_31_n_220 & sub_1130_31_n_22) | ~(sub_1130_31_n_220 | sub_1130_31_n_22));
 assign T_1_11_ = ~((sub_1130_31_n_29 | sub_1130_31_n_28) & ~(sub_1130_31_n_29 & sub_1130_31_n_28));
 assign T_1_20_ = ((sub_1130_31_n_222 & sub_1130_31_n_138) | ~(sub_1130_31_n_222 | sub_1130_31_n_138));
 assign sub_1130_31_n_222 = ~sub_1130_31_n_38;
 assign T_1_32_ = ~(sub_1130_31_n_211 | sub_1130_31_n_193);
 assign sub_1130_31_n_224 = ~(sub_1130_31_n_151 | (sub_1130_31_n_207 & sub_1130_31_n_124));
 assign sub_1130_31_n_223 = ~(sub_1130_31_n_213 & ~sub_1130_31_n_149);
 assign T_1_16_ = ~((sub_1130_31_n_207 | sub_1130_31_n_134) & ~(sub_1130_31_n_207 & sub_1130_31_n_134));
 assign T_1_7_ = ((sub_1130_31_n_209 & sub_1130_31_n_112) | ~(sub_1130_31_n_209 | sub_1130_31_n_112));
 assign T_1_12_ = ~((sub_1130_31_n_39 | sub_1130_31_n_130) & ~(sub_1130_31_n_39 & sub_1130_31_n_130));
 assign T_1_10_ = ((sub_1130_31_n_35 & sub_1130_31_n_16) | ~(sub_1130_31_n_35 | sub_1130_31_n_16));
 assign T_1_9_ = ((sub_1130_31_n_210 & sub_1130_31_n_118) | ~(sub_1130_31_n_210 | sub_1130_31_n_118));
 assign sub_1130_31_n_220 = ~(sub_1130_31_n_57 | (sub_1130_31_n_39 & sub_1130_31_n_70));
 assign sub_1130_31_n_219 = ~(sub_1130_31_n_212 & ~sub_1130_31_n_184);
 assign sub_1130_31_n_213 = ~(sub_1130_31_n_39 & ~sub_1130_31_n_141);
 assign sub_1130_31_n_212 = ~(sub_1130_31_n_208 & ~sub_1130_31_n_169);
 assign sub_1130_31_n_211 = ~(sub_1130_31_n_206 | sub_1130_31_n_182);
 assign sub_1130_31_n_210 = ~(sub_1130_31_n_88 | (~sub_1130_31_n_74 & sub_1130_31_n_198));
 assign sub_1130_31_n_209 = ~(sub_1130_31_n_44 & (~sub_1130_31_n_68 | sub_1130_31_n_199));
 assign sub_1130_31_n_208 = ~sub_1130_31_n_206;
 assign sub_1130_31_n_207 = ~sub_1130_31_n_206;
 assign sub_1130_31_n_206 = ~(sub_1130_31_n_201 | sub_1130_31_n_185);
 assign T_1_6_ = ((sub_1130_31_n_200 & sub_1130_31_n_132) | ~(sub_1130_31_n_200 | sub_1130_31_n_132));
 assign T_1_5_ = ((sub_1130_31_n_196 & sub_1130_31_n_21) | ~(sub_1130_31_n_196 | sub_1130_31_n_21));
 assign T_1_8_ = ~((sub_1130_31_n_198 | sub_1130_31_n_18) & ~(sub_1130_31_n_198 & sub_1130_31_n_18));
 assign sub_1130_31_n_202 = ~(sub_1130_31_n_198 & ~sub_1130_31_n_166);
 assign sub_1130_31_n_201 = ~(sub_1130_31_n_197 | ~sub_1130_31_n_170);
 assign sub_1130_31_n_200 = ~sub_1130_31_n_199;
 assign sub_1130_31_n_199 = ~(sub_1130_31_n_33 | ~sub_1130_31_n_150);
 assign sub_1130_31_n_198 = ~sub_1130_31_n_197;
 assign sub_1130_31_n_197 = ~(sub_1130_31_n_178 | (sub_1130_31_n_190 & sub_1130_31_n_156));
 assign sub_1130_31_n_196 = ~(sub_1130_31_n_100 & (~sub_1130_31_n_3 | sub_1130_31_n_191));
 assign T_1_4_ = ((sub_1130_31_n_191 & sub_1130_31_n_27) | ~(sub_1130_31_n_191 | sub_1130_31_n_27));
 assign T_1_3_ = ~((sub_1130_31_n_189 | sub_1130_31_n_116) & ~(sub_1130_31_n_189 & sub_1130_31_n_116));
 assign sub_1130_31_n_193 = ~(sub_1130_31_n_192 & sub_1130_31_n_187);
 assign sub_1130_31_n_192 = ~(sub_1130_31_n_184 & sub_1130_31_n_174);
 assign sub_1130_31_n_191 = ~sub_1130_31_n_190;
 assign sub_1130_31_n_190 = ~(sub_1130_31_n_186 & sub_1130_31_n_26);
 assign sub_1130_31_n_189 = ~(sub_1130_31_n_14 | (sub_1130_31_n_183 & sub_1130_31_n_67));
 assign T_1_2_ = ~((sub_1130_31_n_183 | sub_1130_31_n_24) & ~(sub_1130_31_n_183 & sub_1130_31_n_24));
 assign sub_1130_31_n_187 = ~(sub_1130_31_n_37 | (sub_1130_31_n_177 & sub_1130_31_n_165));
 assign sub_1130_31_n_186 = ~(sub_1130_31_n_183 & sub_1130_31_n_111);
 assign sub_1130_31_n_185 = ~(sub_1130_31_n_175 & (sub_1130_31_n_180 | sub_1130_31_n_158));
 assign sub_1130_31_n_184 = ~(sub_1130_31_n_176 & (sub_1130_31_n_179 | sub_1130_31_n_159));
 assign sub_1130_31_n_183 = ~(sub_1130_31_n_172 & (sub_1130_31_n_173 & sub_1130_31_n_82));
 assign sub_1130_31_n_182 = ~(sub_1130_31_n_168 & sub_1130_31_n_174);
 assign T_1_1_ = ~((sub_1130_31_n_113 | n_1359) & ~(sub_1130_31_n_113 & n_1359));
 assign sub_1130_31_n_180 = ~(sub_1130_31_n_157 | (sub_1130_31_n_153 & sub_1130_31_n_136));
 assign sub_1130_31_n_179 = ~(sub_1130_31_n_145 | (sub_1130_31_n_151 & sub_1130_31_n_128));
 assign sub_1130_31_n_178 = ~(sub_1130_31_n_154 & (sub_1130_31_n_150 | sub_1130_31_n_121));
 assign sub_1130_31_n_177 = ~(sub_1130_31_n_171 & ~sub_1130_31_n_147);
 assign sub_1130_31_n_176 = ~(sub_1130_31_n_144 | (sub_1130_31_n_160 & sub_1130_31_n_143));
 assign sub_1130_31_n_175 = ~(sub_1130_31_n_146 | (sub_1130_31_n_149 & sub_1130_31_n_117));
 assign sub_1130_31_n_174 = ~(sub_1130_31_n_162 | sub_1130_31_n_164);
 assign sub_1130_31_n_173 = ~(n_1359 & R_2_0_);
 assign sub_1130_31_n_172 = ~(n_1359 & ~n_1353);
 assign sub_1130_31_n_171 = ~(sub_1130_31_n_152 & ~sub_1130_31_n_137);
 assign sub_1130_31_n_170 = ~(sub_1130_31_n_166 | sub_1130_31_n_158);
 assign sub_1130_31_n_169 = ~sub_1130_31_n_168;
 assign sub_1130_31_n_168 = ~(sub_1130_31_n_161 | sub_1130_31_n_159);
 assign sub_1130_31_n_167 = ~(sub_1130_31_n_148 & sub_1130_31_n_122);
 assign sub_1130_31_n_165 = ~sub_1130_31_n_164;
 assign sub_1130_31_n_163 = ~sub_1130_31_n_162;
 assign sub_1130_31_n_157 = ~(sub_1130_31_n_8 & (sub_1130_31_n_55 | sub_1130_31_n_94));
 assign sub_1130_31_n_156 = ~(sub_1130_31_n_120 | sub_1130_31_n_121);
 assign sub_1130_31_n_155 = ~(sub_1130_31_n_32 & sub_1130_31_n_54);
 assign sub_1130_31_n_154 = ~(sub_1130_31_n_105 | (sub_1130_31_n_86 & sub_1130_31_n_12));
 assign sub_1130_31_n_166 = ~(sub_1130_31_n_139 & sub_1130_31_n_136);
 assign sub_1130_31_n_164 = ~(sub_1130_31_n_126 & sub_1130_31_n_0);
 assign sub_1130_31_n_162 = ~(sub_1130_31_n_125 & ~sub_1130_31_n_137);
 assign sub_1130_31_n_161 = ~(sub_1130_31_n_124 & sub_1130_31_n_128);
 assign sub_1130_31_n_160 = ~(sub_1130_31_n_104 & (sub_1130_31_n_101 | sub_1130_31_n_87));
 assign sub_1130_31_n_159 = ~(sub_1130_31_n_142 & sub_1130_31_n_143);
 assign sub_1130_31_n_158 = ~(sub_1130_31_n_140 & sub_1130_31_n_117);
 assign sub_1130_31_n_147 = ~(sub_1130_31_n_80 & (sub_1130_31_n_89 | sub_1130_31_n_91));
 assign sub_1130_31_n_146 = ~(sub_1130_31_n_81 & (sub_1130_31_n_10 | sub_1130_31_n_93));
 assign sub_1130_31_n_145 = ~(sub_1130_31_n_106 & (sub_1130_31_n_98 | sub_1130_31_n_63));
 assign sub_1130_31_n_144 = ~(sub_1130_31_n_108 & (sub_1130_31_n_54 | sub_1130_31_n_95));
 assign sub_1130_31_n_153 = ~(sub_1130_31_n_5 & (sub_1130_31_n_13 | sub_1130_31_n_96));
 assign sub_1130_31_n_152 = ~(sub_1130_31_n_4 & (~sub_1130_31_n_71 | sub_1130_31_n_58));
 assign sub_1130_31_n_151 = ~(sub_1130_31_n_11 & (sub_1130_31_n_76 | sub_1130_31_n_77));
 assign sub_1130_31_n_150 = ~(sub_1130_31_n_78 | (sub_1130_31_n_99 & sub_1130_31_n_6));
 assign sub_1130_31_n_149 = ~(sub_1130_31_n_83 & (sub_1130_31_n_56 | sub_1130_31_n_61));
 assign sub_1130_31_n_148 = ~(sub_1130_31_n_110 | ~sub_1130_31_n_79);
 assign sub_1130_31_n_141 = ~sub_1130_31_n_140;
 assign sub_1130_31_n_129 = ~(sub_1130_31_n_9 & ~n_1276);
 assign sub_1130_31_n_143 = ~(sub_1130_31_n_97 | sub_1130_31_n_95);
 assign sub_1130_31_n_142 = ~(sub_1130_31_n_59 | sub_1130_31_n_87);
 assign sub_1130_31_n_140 = ~(sub_1130_31_n_69 | sub_1130_31_n_61);
 assign sub_1130_31_n_139 = ~(sub_1130_31_n_74 | sub_1130_31_n_96);
 assign sub_1130_31_n_138 = (sub_1130_31_n_101 & sub_1130_31_n_60);
 assign sub_1130_31_n_137 = ~(sub_1130_31_n_15 & sub_1130_31_n_92);
 assign sub_1130_31_n_136 = ~(sub_1130_31_n_45 | sub_1130_31_n_94);
 assign sub_1130_31_n_135 = (sub_1130_31_n_98 & sub_1130_31_n_85);
 assign sub_1130_31_n_134 = ~(sub_1130_31_n_76 & sub_1130_31_n_103);
 assign sub_1130_31_n_133 = ~(sub_1130_31_n_93 | ~sub_1130_31_n_81);
 assign sub_1130_31_n_132 = ~(sub_1130_31_n_44 & sub_1130_31_n_68);
 assign sub_1130_31_n_131 = ~(sub_1130_31_n_10 & sub_1130_31_n_65);
 assign sub_1130_31_n_130 = ~(sub_1130_31_n_56 & sub_1130_31_n_70);
 assign sub_1130_31_n_123 = ~sub_1130_31_n_122;
 assign sub_1130_31_n_111 = ~(sub_1130_31_n_66 | sub_1130_31_n_90);
 assign sub_1130_31_n_110 = ~(sub_1130_31_n_1 | ~sub_1130_31_n_2);
 assign T_1_0_ = ~(sub_1130_31_n_53 & (~{in2[1]} | {in1[0]}));
 assign sub_1130_31_n_128 = ~(sub_1130_31_n_84 | sub_1130_31_n_63);
 assign sub_1130_31_n_127 = ~(sub_1130_31_n_79 & sub_1130_31_n_2);
 assign sub_1130_31_n_126 = ~(sub_1130_31_n_75 | ~sub_1130_31_n_2);
 assign sub_1130_31_n_125 = ~(sub_1130_31_n_72 | ~sub_1130_31_n_71);
 assign sub_1130_31_n_124 = ~(sub_1130_31_n_102 | sub_1130_31_n_77);
 assign sub_1130_31_n_122 = ~(sub_1130_31_n_9 | sub_1130_31_n_107);
 assign sub_1130_31_n_121 = ~(sub_1130_31_n_68 & sub_1130_31_n_12);
 assign sub_1130_31_n_120 = ~(sub_1130_31_n_3 & sub_1130_31_n_6);
 assign sub_1130_31_n_119 = ~(sub_1130_31_n_80 & sub_1130_31_n_92);
 assign sub_1130_31_n_118 = ~(sub_1130_31_n_96 | ~sub_1130_31_n_5);
 assign sub_1130_31_n_117 = ~(sub_1130_31_n_64 | sub_1130_31_n_93);
 assign sub_1130_31_n_116 = ~(sub_1130_31_n_43 | sub_1130_31_n_90);
 assign sub_1130_31_n_115 = ~(sub_1130_31_n_4 & sub_1130_31_n_71);
 assign sub_1130_31_n_114 = ~(sub_1130_31_n_58 & sub_1130_31_n_73);
 assign sub_1130_31_n_113 = ~(sub_1130_31_n_82 & sub_1130_31_n_7);
 assign sub_1130_31_n_112 = ~(sub_1130_31_n_46 & sub_1130_31_n_12);
 assign sub_1130_31_n_105 = ~sub_1130_31_n_46;
 assign sub_1130_31_n_103 = ~sub_1130_31_n_102;
 assign sub_1130_31_n_100 = ~sub_1130_31_n_99;
 assign sub_1130_31_n_92 = ~sub_1130_31_n_91;
 assign sub_1130_31_n_88 = ~sub_1130_31_n_13;
 assign sub_1130_31_n_86 = ~sub_1130_31_n_44;
 assign sub_1130_31_n_85 = ~sub_1130_31_n_84;
 assign sub_1130_31_n_108 = ~(R_2_22_ & ~n_1295);
 assign sub_1130_31_n_107 = ~(R_2_29_ | ~n_833);
 assign sub_1130_31_n_106 = ~(R_2_18_ & ~n_1305);
 assign sub_1130_31_n_46 = ~(R_2_6_ & ~n_1170);
 assign sub_1130_31_n_104 = ~(R_2_20_ & ~n_1369);
 assign sub_1130_31_n_102 = ~(R_2_15_ | ~n_1139);
 assign sub_1130_31_n_101 = ~(R_2_19_ & ~n_1215);
 assign sub_1130_31_n_99 = ~(n_1343 | sub_1130_31_n_52);
 assign sub_1130_31_n_98 = ~(R_2_17_ & ~n_1034);
 assign sub_1130_31_n_97 = ~(R_2_21_ | ~n_1180);
 assign sub_1130_31_n_96 = ~(R_2_8_ | ~n_1165);
 assign sub_1130_31_n_45 = ~(R_2_9_ | ~n_1348);
 assign sub_1130_31_n_95 = ~(R_2_22_ | ~n_1295);
 assign sub_1130_31_n_94 = ~(R_2_10_ | ~n_1068);
 assign sub_1130_31_n_93 = ~(R_2_14_ | ~n_1094);
 assign sub_1130_31_n_91 = ~(R_2_26_ | ~n_1245);
 assign sub_1130_31_n_90 = ~(R_2_2_ | ~n_1116);
 assign sub_1130_31_n_89 = ~(R_2_25_ & ~n_1089);
 assign sub_1130_31_n_87 = ~(R_2_20_ | ~n_1369);
 assign sub_1130_31_n_44 = ~(sub_1130_31_n_51 & R_2_5_);
 assign sub_1130_31_n_84 = ~(R_2_17_ | ~n_1034);
 assign sub_1130_31_n_73 = ~sub_1130_31_n_72;
 assign sub_1130_31_n_70 = ~sub_1130_31_n_69;
 assign sub_1130_31_n_67 = ~sub_1130_31_n_66;
 assign sub_1130_31_n_65 = ~sub_1130_31_n_64;
 assign sub_1130_31_n_62 = ~sub_1130_31_n_10;
 assign sub_1130_31_n_60 = ~sub_1130_31_n_59;
 assign sub_1130_31_n_57 = ~sub_1130_31_n_56;
 assign sub_1130_31_n_83 = ~(R_2_12_ & ~n_1262);
 assign sub_1130_31_n_82 = ~(R_2_0_ & ~n_1353);
 assign sub_1130_31_n_81 = ~(R_2_14_ & ~n_1094);
 assign sub_1130_31_n_80 = ~(R_2_26_ & ~n_1245);
 assign sub_1130_31_n_79 = ~(sub_1130_31_n_48 & R_2_28_);
 assign sub_1130_31_n_78 = ~(n_1052 | sub_1130_31_n_47);
 assign sub_1130_31_n_77 = ~(R_2_16_ | ~n_1175);
 assign sub_1130_31_n_76 = ~(R_2_15_ & ~n_1139);
 assign sub_1130_31_n_75 = ~(R_2_27_ | ~n_1300);
 assign sub_1130_31_n_74 = ~(R_2_7_ | ~n_1220);
 assign sub_1130_31_n_72 = ~(R_2_23_ | ~n_1062);
 assign sub_1130_31_n_71 = ~(sub_1130_31_n_50 & n_1374);
 assign sub_1130_31_n_69 = ~(R_2_11_ | ~n_1029);
 assign sub_1130_31_n_68 = ~(sub_1130_31_n_49 & ~sub_1130_31_n_51);
 assign sub_1130_31_n_66 = ~(R_2_1_ | ~n_1104);
 assign sub_1130_31_n_64 = ~(R_2_13_ | ~n_1185);
 assign sub_1130_31_n_63 = ~(R_2_18_ | ~n_1305);
 assign sub_1130_31_n_61 = ~(R_2_12_ | ~n_1262);
 assign sub_1130_31_n_59 = ~(R_2_19_ | ~n_1215);
 assign sub_1130_31_n_58 = ~(R_2_23_ & ~n_1062);
 assign sub_1130_31_n_56 = ~(R_2_11_ & ~n_1029);
 assign sub_1130_31_n_55 = ~(R_2_9_ & ~n_1348);
 assign sub_1130_31_n_54 = ~(R_2_21_ & ~n_1180);
 assign sub_1130_31_n_53 = ~({in1[0]} & ~{in2[1]});
 assign sub_1130_31_n_52 = ~R_2_3_;
 assign sub_1130_31_n_51 = ~n_1099;
 assign sub_1130_31_n_50 = ~R_2_24_;
 assign sub_1130_31_n_49 = ~R_2_5_;
 assign sub_1130_31_n_48 = ~n_1364;
 assign sub_1130_31_n_47 = ~R_2_4_;
 assign sub_1130_31_n_43 = ~(n_1116 | ~R_2_2_);
 assign sub_1130_31_n_42 = (sub_1130_31_n_32 | (sub_1130_31_n_54 & sub_1130_31_n_239));
 assign sub_1130_31_n_41 = ~(sub_1130_31_n_58 & ~(sub_1130_31_n_73 & sub_1130_31_n_219));
 assign sub_1130_31_n_40 = ~(sub_1130_31_n_76 & ~(sub_1130_31_n_103 & sub_1130_31_n_207));
 assign sub_1130_31_n_39 = ~(sub_1130_31_n_202 & sub_1130_31_n_180);
 assign sub_1130_31_n_38 = ~(sub_1130_31_n_179 & (sub_1130_31_n_161 | sub_1130_31_n_206));
 assign sub_1130_31_n_37 = ~(sub_1130_31_n_129 & (~sub_1130_31_n_0 | sub_1130_31_n_148));
 assign sub_1130_31_n_36 = ~(sub_1130_31_n_38 & sub_1130_31_n_142);
 assign sub_1130_31_n_35 = ~(sub_1130_31_n_153 | (sub_1130_31_n_139 & sub_1130_31_n_198));
 assign sub_1130_31_n_34 = ~(sub_1130_31_n_152 | (sub_1130_31_n_125 & sub_1130_31_n_219));
 assign sub_1130_31_n_33 = ~(sub_1130_31_n_191 | sub_1130_31_n_120);
 assign sub_1130_31_n_32 = ~(sub_1130_31_n_95 | ~sub_1130_31_n_108);
 assign sub_1130_31_n_31 = ~(sub_1130_31_n_75 | ~sub_1130_31_n_1);
 assign sub_1130_31_n_30 = ~(sub_1130_31_n_54 & ~sub_1130_31_n_97);
 assign sub_1130_31_n_29 = ~(sub_1130_31_n_55 & (sub_1130_31_n_45 | sub_1130_31_n_35));
 assign sub_1130_31_n_28 = ~(sub_1130_31_n_8 & ~sub_1130_31_n_94);
 assign sub_1130_31_n_27 = ~(sub_1130_31_n_99 | ~sub_1130_31_n_3);
 assign sub_1130_31_n_26 = ~(sub_1130_31_n_43 | (~sub_1130_31_n_90 & sub_1130_31_n_14));
 assign sub_1130_31_n_25 = (sub_1130_31_n_89 & sub_1130_31_n_15);
 assign sub_1130_31_n_24 = ~(sub_1130_31_n_67 & ~sub_1130_31_n_14);
 assign sub_1130_31_n_23 = ~(sub_1130_31_n_104 & ~sub_1130_31_n_87);
 assign sub_1130_31_n_22 = ~(sub_1130_31_n_61 | ~sub_1130_31_n_83);
 assign sub_1130_31_n_21 = ~(sub_1130_31_n_6 & ~sub_1130_31_n_78);
 assign sub_1130_31_n_20 = ~(sub_1130_31_n_11 & ~sub_1130_31_n_77);
 assign sub_1130_31_n_19 = ~(sub_1130_31_n_1 & (sub_1130_31_n_75 | sub_1130_31_n_232));
 assign sub_1130_31_n_18 = ~(sub_1130_31_n_13 & ~sub_1130_31_n_74);
 assign sub_1130_31_n_17 = ~(sub_1130_31_n_106 & ~sub_1130_31_n_63);
 assign sub_1130_31_n_16 = ~(sub_1130_31_n_45 | ~sub_1130_31_n_55);
 assign sub_1130_31_n_15 = ~(n_1089 & ~R_2_25_);
 assign sub_1130_31_n_14 = ~(n_1104 | ~R_2_1_);
 assign sub_1130_31_n_13 = ~(R_2_7_ & ~n_1220);
 assign sub_1130_31_n_12 = ~(n_1170 & ~R_2_6_);
 assign sub_1130_31_n_11 = ~(R_2_16_ & ~n_1175);
 assign sub_1130_31_n_10 = ~(R_2_13_ & ~n_1185);
 assign sub_1130_31_n_9 = ~(n_833 | ~R_2_29_);
 assign sub_1130_31_n_8 = ~(R_2_10_ & ~n_1068);
 assign sub_1130_31_n_7 = ~(n_1353 & ~R_2_0_);
 assign sub_1130_31_n_6 = ~(sub_1130_31_n_47 & n_1052);
 assign sub_1130_31_n_5 = ~(R_2_8_ & ~n_1165);
 assign sub_1130_31_n_4 = (sub_1130_31_n_50 | n_1374);
 assign sub_1130_31_n_3 = ~(sub_1130_31_n_52 & n_1343);
 assign sub_1130_31_n_2 = (R_2_28_ | sub_1130_31_n_48);
 assign sub_1130_31_n_1 = ~(R_2_27_ & ~n_1300);
 assign sub_1130_31_n_0 = ~(sub_1130_31_n_107 | n_1276);
 assign T_0_32_ = ~(sub_1160_30_n_122 | (sub_1160_30_n_123 | sub_1160_30_n_125));
 assign sub_1160_30_n_125 = ~(sub_1160_30_n_124 | (sub_1160_30_n_114 | sub_1160_30_n_108));
 assign sub_1160_30_n_124 = ~(sub_1160_30_n_119 | (sub_1160_30_n_107 & (sub_1160_30_n_79 & sub_1160_30_n_121)));
 assign sub_1160_30_n_123 = ~(sub_1160_30_n_116 & (sub_1160_30_n_98 & sub_1160_30_n_118));
 assign sub_1160_30_n_122 = ~(sub_1160_30_n_114 | sub_1160_30_n_120);
 assign sub_1160_30_n_121 = ~(sub_1160_30_n_112 & (sub_1160_30_n_86 | sub_1160_30_n_115));
 assign sub_1160_30_n_120 = ~(sub_1160_30_n_109 | (sub_1160_30_n_111 & sub_1160_30_n_95));
 assign sub_1160_30_n_119 = ~(sub_1160_30_n_110 & (sub_1160_30_n_113 | sub_1160_30_n_94));
 assign sub_1160_30_n_118 = ~(sub_1160_30_n_81 & (sub_1160_30_n_74 & sub_1160_30_n_117));
 assign sub_1160_30_n_117 = ~(sub_1160_30_n_102 & (sub_1160_30_n_105 | sub_1160_30_n_76));
 assign sub_1160_30_n_116 = ~(sub_1160_30_n_74 & ~sub_1160_30_n_106);
 assign sub_1160_30_n_115 = ~(sub_1160_30_n_92 | (sub_1160_30_n_88 & sub_1160_30_n_70));
 assign sub_1160_30_n_114 = ~(sub_1160_30_n_87 & (sub_1160_30_n_96 & sub_1160_30_n_74));
 assign sub_1160_30_n_113 = ~(sub_1160_30_n_100 | (sub_1160_30_n_99 & sub_1160_30_n_85));
 assign sub_1160_30_n_112 = ~(sub_1160_30_n_97 | (sub_1160_30_n_93 & sub_1160_30_n_77));
 assign sub_1160_30_n_111 = ~(sub_1160_30_n_104 & (sub_1160_30_n_91 | sub_1160_30_n_75));
 assign sub_1160_30_n_110 = ~(sub_1160_30_n_90 | (sub_1160_30_n_103 & sub_1160_30_n_83));
 assign sub_1160_30_n_109 = ~(sub_1160_30_n_89 & (sub_1160_30_n_101 | sub_1160_30_n_84));
 assign sub_1160_30_n_108 = ~(sub_1160_30_n_95 & (sub_1160_30_n_4 & ~sub_1160_30_n_75));
 assign sub_1160_30_n_107 = ~(sub_1160_30_n_94 | ~sub_1160_30_n_85);
 assign sub_1160_30_n_106 = ~((sub_1160_30_n_19 & R_1_28_) | (R_1_27_ & sub_1160_30_n_73));
 assign sub_1160_30_n_105 = ~((sub_1160_30_n_30 & R_1_24_) | (sub_1160_30_n_78 & R_1_23_));
 assign sub_1160_30_n_104 = ~((sub_1160_30_n_8 & R_1_18_) | (sub_1160_30_n_36 & sub_1160_30_n_3));
 assign sub_1160_30_n_103 = ~((n_1262 | sub_1160_30_n_7) & (sub_1160_30_n_33 | sub_1160_30_n_45));
 assign sub_1160_30_n_102 = ~((sub_1160_30_n_31 & R_1_26_) | (sub_1160_30_n_61 & sub_1160_30_n_57));
 assign sub_1160_30_n_101 = ~(sub_1160_30_n_50 | (sub_1160_30_n_26 & (R_1_19_ & sub_1160_30_n_65)));
 assign sub_1160_30_n_100 = ~((n_1068 | sub_1160_30_n_9) & (sub_1160_30_n_38 | sub_1160_30_n_66));
 assign sub_1160_30_n_99 = ~((n_1165 | sub_1160_30_n_28) & (sub_1160_30_n_34 | sub_1160_30_n_64));
 assign sub_1160_30_n_98 = ~((sub_1160_30_n_13 & R_1_30_) | (sub_1160_30_n_2 & sub_1160_30_n_47));
 assign sub_1160_30_n_97 = ~((n_1170 | sub_1160_30_n_21) & (sub_1160_30_n_51 | sub_1160_30_n_49));
 assign sub_1160_30_n_96 = ~(sub_1160_30_n_76 | (sub_1160_30_n_15 & n_1062));
 assign sub_1160_30_n_93 = ~((n_1052 | sub_1160_30_n_24) & (sub_1160_30_n_60 | sub_1160_30_n_68));
 assign sub_1160_30_n_92 = ~((n_1116 | sub_1160_30_n_14) & (sub_1160_30_n_0 | sub_1160_30_n_41));
 assign sub_1160_30_n_91 = ~(sub_1160_30_n_1 | (sub_1160_30_n_20 & (R_1_15_ & sub_1160_30_n_48)));
 assign sub_1160_30_n_90 = ~((n_1094 | sub_1160_30_n_17) & (sub_1160_30_n_58 | sub_1160_30_n_42));
 assign sub_1160_30_n_89 = ~((sub_1160_30_n_32 & R_1_22_) | (sub_1160_30_n_67 & sub_1160_30_n_69));
 assign sub_1160_30_n_88 = ~((n_1281 & sub_1160_30_n_16) | ((sub_1160_30_n_16 & n_1353) | (n_1353 & n_1281)));
 assign sub_1160_30_n_87 = ~(sub_1160_30_n_80 | sub_1160_30_n_43);
 assign sub_1160_30_n_86 = ~(sub_1160_30_n_71 & sub_1160_30_n_77);
 assign sub_1160_30_n_95 = ~(sub_1160_30_n_72 | sub_1160_30_n_84);
 assign sub_1160_30_n_94 = ~(sub_1160_30_n_82 & sub_1160_30_n_83);
 assign sub_1160_30_n_82 = ~(sub_1160_30_n_53 | sub_1160_30_n_45);
 assign sub_1160_30_n_81 = ~(sub_1160_30_n_43 | ~sub_1160_30_n_44);
 assign sub_1160_30_n_80 = ~(sub_1160_30_n_63 & sub_1160_30_n_44);
 assign sub_1160_30_n_79 = ~(sub_1160_30_n_37 | sub_1160_30_n_64);
 assign sub_1160_30_n_78 = ~(sub_1160_30_n_62 | n_1062);
 assign sub_1160_30_n_85 = ~(sub_1160_30_n_66 | (sub_1160_30_n_6 & n_1348));
 assign sub_1160_30_n_84 = ~(sub_1160_30_n_67 & (R_1_21_ | sub_1160_30_n_12));
 assign sub_1160_30_n_83 = ~(sub_1160_30_n_59 | sub_1160_30_n_42);
 assign sub_1160_30_n_73 = ~(sub_1160_30_n_39 & (n_1300 | n_1364));
 assign sub_1160_30_n_72 = ~(sub_1160_30_n_65 & (R_1_19_ | sub_1160_30_n_26));
 assign sub_1160_30_n_71 = ~(sub_1160_30_n_35 | sub_1160_30_n_68);
 assign sub_1160_30_n_70 = ~(sub_1160_30_n_40 | sub_1160_30_n_41);
 assign sub_1160_30_n_77 = ~(sub_1160_30_n_49 | (~R_1_5_ & ~sub_1160_30_n_22));
 assign sub_1160_30_n_76 = ~(sub_1160_30_n_61 & (R_1_25_ | sub_1160_30_n_11));
 assign sub_1160_30_n_75 = ~(sub_1160_30_n_52 & sub_1160_30_n_3);
 assign sub_1160_30_n_74 = ~(sub_1160_30_n_54 | sub_1160_30_n_46);
 assign sub_1160_30_n_69 = ~sub_1160_30_n_55;
 assign sub_1160_30_n_63 = ~sub_1160_30_n_62;
 assign sub_1160_30_n_60 = ~(R_1_3_ & ~n_1343);
 assign sub_1160_30_n_59 = ~(R_1_13_ | ~n_1185);
 assign sub_1160_30_n_58 = ~(R_1_13_ & ~n_1185);
 assign sub_1160_30_n_57 = (sub_1160_30_n_11 & R_1_25_);
 assign sub_1160_30_n_56 = ~({in2[0]} | ~{in1[0]});
 assign sub_1160_30_n_55 = ~(sub_1160_30_n_12 & R_1_21_);
 assign sub_1160_30_n_54 = ~(R_1_29_ | ~n_833);
 assign sub_1160_30_n_53 = ~(R_1_11_ | ~n_1029);
 assign sub_1160_30_n_52 = ~(sub_1160_30_n_23 & n_1034);
 assign sub_1160_30_n_51 = ~(sub_1160_30_n_22 & R_1_5_);
 assign sub_1160_30_n_50 = ~(n_1369 | sub_1160_30_n_27);
 assign sub_1160_30_n_68 = ~(R_1_4_ | ~n_1052);
 assign sub_1160_30_n_67 = ~(sub_1160_30_n_10 & ~sub_1160_30_n_32);
 assign sub_1160_30_n_66 = ~(R_1_10_ | ~n_1068);
 assign sub_1160_30_n_65 = ~(sub_1160_30_n_27 & n_1369);
 assign sub_1160_30_n_64 = ~(R_1_8_ | ~n_1165);
 assign sub_1160_30_n_62 = ~(R_1_24_ | ~n_1374);
 assign sub_1160_30_n_61 = ~(sub_1160_30_n_29 & ~sub_1160_30_n_31);
 assign sub_1160_30_n_47 = ~sub_1160_30_n_46;
 assign sub_1160_30_n_40 = ~(R_1_1_ | ~n_1104);
 assign sub_1160_30_n_39 = ~(R_1_28_ & ~n_1300);
 assign sub_1160_30_n_38 = ~(R_1_9_ & ~n_1348);
 assign sub_1160_30_n_37 = ~(R_1_7_ | ~n_1220);
 assign sub_1160_30_n_36 = ~(n_1034 | sub_1160_30_n_23);
 assign sub_1160_30_n_35 = ~(R_1_3_ | ~n_1343);
 assign sub_1160_30_n_34 = ~(sub_1160_30_n_25 & R_1_7_);
 assign sub_1160_30_n_33 = ~(R_1_11_ & ~n_1029);
 assign sub_1160_30_n_49 = ~(R_1_6_ | ~n_1170);
 assign sub_1160_30_n_48 = ~(n_1175 & ~R_1_16_);
 assign sub_1160_30_n_46 = ~(R_1_30_ | ~n_1276);
 assign sub_1160_30_n_45 = ~(R_1_12_ | ~n_1262);
 assign sub_1160_30_n_44 = ~(sub_1160_30_n_18 & ~sub_1160_30_n_19);
 assign sub_1160_30_n_43 = ~(R_1_27_ | ~n_1300);
 assign sub_1160_30_n_42 = ~(R_1_14_ | ~n_1094);
 assign sub_1160_30_n_41 = ~(R_1_2_ | ~n_1116);
 assign sub_1160_30_n_32 = ~n_1295;
 assign sub_1160_30_n_31 = ~n_1245;
 assign sub_1160_30_n_30 = ~n_1374;
 assign sub_1160_30_n_29 = ~R_1_26_;
 assign sub_1160_30_n_28 = ~R_1_8_;
 assign sub_1160_30_n_27 = ~R_1_20_;
 assign sub_1160_30_n_26 = ~n_1215;
 assign sub_1160_30_n_25 = ~n_1220;
 assign sub_1160_30_n_24 = ~R_1_4_;
 assign sub_1160_30_n_23 = ~R_1_17_;
 assign sub_1160_30_n_22 = ~n_1099;
 assign sub_1160_30_n_21 = ~R_1_6_;
 assign sub_1160_30_n_20 = ~n_1139;
 assign sub_1160_30_n_19 = ~n_1364;
 assign sub_1160_30_n_18 = ~R_1_28_;
 assign sub_1160_30_n_17 = ~R_1_14_;
 assign sub_1160_30_n_16 = ~R_1_0_;
 assign sub_1160_30_n_15 = ~R_1_23_;
 assign sub_1160_30_n_14 = ~R_1_2_;
 assign sub_1160_30_n_13 = ~n_1276;
 assign sub_1160_30_n_12 = ~n_1180;
 assign sub_1160_30_n_11 = ~n_1089;
 assign sub_1160_30_n_10 = ~R_1_22_;
 assign sub_1160_30_n_9 = ~R_1_10_;
 assign sub_1160_30_n_8 = ~n_1305;
 assign sub_1160_30_n_7 = ~R_1_12_;
 assign sub_1160_30_n_6 = ~R_1_9_;
 assign sub_1160_30_n_4 = (sub_1160_30_n_48 & (R_1_15_ | sub_1160_30_n_20));
 assign sub_1160_30_n_3 = (R_1_18_ | sub_1160_30_n_8);
 assign sub_1160_30_n_2 = ~(n_833 | ~R_1_29_);
 assign sub_1160_30_n_1 = ~(n_1175 | ~R_1_16_);
 assign sub_1160_30_n_0 = ~(R_1_1_ & ~n_1104);
endmodule



